.SUBCKT INVD1 I ZN
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.96e-07  AD=6.4e-14  AS=8.4e-14  PD=1.11e-06  PS=1.21e-06  SA=2.15e-07  SB=1.65e-07  NRD=0.474  NRS=0.668  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vdd vdd pch L=6e-08 W=5.23e-07  AD=8.6e-14  AS=1.12e-13  PD=1.37e-06  PS=1.47e-06  SA=2.15e-07  SB=1.65e-07  NRD=0.433  NRS=0.58  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M1:DRN ZN 15.2446 
CC38171 M1:DRN M1:GATE 3.864e-17
CC38168 M1:DRN I 8.83e-18
R1 ZN M2:DRN 15.3531 
CC38170 ZN M1:GATE 1.03e-18
CC38165 ZN M2:GATE 1.085e-17
CC38169 ZN I 3.149e-17
CC38166 M2:DRN M2:GATE 4.32e-17
CC38167 M2:DRN I 4.85e-18
C2 M1:DRN 0 2.382e-17
C3 ZN 0 1.4107e-16
C4 M2:DRN 0 2.864e-17
R5 M2:GATE I 200.165 
R6 I M1:GATE 169.187 
R7 M1:GATE M2:GATE 462.598 
C8 I 0 1.1015e-16
C9 M1:GATE 0 4.87e-17
C10 M2:GATE 0 9.383e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
