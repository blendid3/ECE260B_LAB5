.SUBCKT NR2D4 A1 A2 ZN
MMM10 M9:SRC M10:GATE M10:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.75e-06  SB=4.5e-07  NRD=2.009  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 M11:DRN M11:GATE M11:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.49e-06  SB=7.1e-07  NRD=2.099  NRS=2.009  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7.4e-14  AS=3.9e-14  PD=1.16e-06  PS=5.9e-07  SA=2.015e-06  SB=1.9e-07  NRD=0.619  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M11:SRC M12:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.23e-06  SB=9.7e-07  NRD=2.009  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.745e-06  SB=4.5e-07  NRD=4.183  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=9.9e-07  SB=1.21e-06  NRD=6.61  NRS=2.009  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.485e-06  SB=7.1e-07  NRD=4.537  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M13:SRC M14:GATE M14:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7.3e-07  SB=1.47e-06  NRD=2.009  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=1.225e-06  SB=9.7e-07  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 M15:DRN M15:GATE M15:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.7e-07  SB=1.73e-06  NRD=2.099  NRS=2.009  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=9.85e-07  SB=1.21e-06  NRD=7.648  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M15:SRC M16:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=1.09e-13  PD=7.2e-07  PS=1.46e-06  SA=2.1e-07  SB=1.99e-06  NRD=2.009  NRS=0.495  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.25e-07  SB=1.47e-06  NRD=4.183  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.65e-07  SB=1.73e-06  NRD=4.537  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=8e-14  PD=5.9e-07  PS=1.19e-06  SA=2.05e-07  SB=1.99e-06  NRD=4.183  NRS=0.566  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.2e-07  AD=9.9e-14  AS=5.2e-14  PD=1.42e-06  PS=7.2e-07  SA=2.01e-06  SB=1.9e-07  NRD=0.466  NRS=2.009  SCA=9.643  SCB=0.01  SCC=0.000823 
CC47812 M9:SRC A2:1 1.08e-18
R0 ZN:2 M5:SRC 79.1107 
R1 ZN:1 M5:SRC 49.2604 
R2 M5:SRC M6:DRN 0.001 
CC47877 M5:SRC M5:GATE 4.57e-18
CC47798 M5:SRC M6:GATE 4.57e-18
CC47782 M5:SRC A1 1.571e-17
CC47830 M5:SRC A2:2 2.646e-17
CC47757 M5:SRC A1:1 1.714e-17
R3 M7:SRC ZN:1 29.9999 
R4 M3:SRC ZN:1 127.35 
R5 ZN:2 ZN:1 1.103 
R6 ZN:1 M14:SRC 31.5109 
CC47795 ZN:1 M3:GATE 1.9e-18
CC47799 ZN:1 M6:GATE 7.53e-18
CC47790 ZN:1 M2:GATE 5.17e-18
CC47881 ZN:1 M5:GATE 1.93e-18
CC47889 ZN:1 M4:GATE 1.93e-18
CC47785 ZN:1 A1 7.424e-17
CC47857 ZN:1 M12:GATE 3.79e-18
CC47835 ZN:1 A2:2 3.26e-18
CC47842 ZN:1 M16:GATE 3.34e-18
CC47803 ZN:1 M7:GATE 2.09e-18
CC47819 ZN:1 A2:1 1.2e-16
CC47758 ZN:1 A1:1 1.331e-17
CC47905 ZN:1 M1:GATE 3.75e-18
CC47771 ZN:1 M14:GATE 3.6e-18
CC47766 ZN:1 A1:2 2.88e-18
CC47769 ZN:1 M15:GATE 8.78e-18
CC47896 ZN:1 M8:GATE 6.92e-18
R7 M14:SRC M15:DRN 0.001 
CC47807 M14:SRC A2:1 1.061e-17
CC47755 M14:SRC A1:1 9.48e-18
CC47779 M14:SRC A1 3.25e-18
CC47768 M14:SRC M15:GATE 2.78e-17
CC47770 M14:SRC M14:GATE 2.82e-17
R8 M1:SRC ZN:2 30.0801 
R9 ZN ZN:2 0.09797 
R10 ZN:2 M3:SRC 39.5835 
CC47796 ZN:2 M3:GATE 1.48e-18
CC47786 ZN:2 A1 7.926e-17
CC47791 ZN:2 M2:GATE 1.62e-18
CC47838 ZN:2 A2:2 4.48e-18
CC47804 ZN:2 M7:GATE 1.43e-18
CC47759 ZN:2 A1:1 2.4e-18
CC47891 ZN:2 M4:GATE 1.12e-18
CC47767 ZN:2 A1:2 3.01e-18
CC47898 ZN:2 M8:GATE 3.46e-18
R11 M3:SRC M4:DRN 0.001 
CC47885 M3:SRC M4:GATE 4.57e-18
CC47792 M3:SRC M3:GATE 4.57e-18
CC47783 M3:SRC A1 3.08e-18
CC47831 M3:SRC A2:2 2.443e-17
CC47763 M3:SRC A1:2 2.653e-17
R12 ZN M10:SRC 30.8024 
R13 M10:SRC M11:DRN 0.001 
CC47810 M10:SRC A2:1 4.87e-18
CC47762 M10:SRC A1:2 1.142e-17
CC47774 M10:SRC M11:GATE 2.801e-17
CC47777 M10:SRC M10:GATE 2.769e-17
CC47789 ZN M2:GATE 5.45e-18
CC47784 ZN A1 5.167e-17
CC47794 ZN M3:GATE 2.26e-18
CC47833 ZN A2:2 1.04e-18
CC47855 ZN M12:GATE 1.03e-18
CC47865 ZN M9:GATE 1.68e-18
CC47817 ZN A2:1 9.711e-17
CC47903 ZN M1:GATE 3.28e-18
CC47775 ZN M11:GATE 7.43e-18
CC47778 ZN M10:GATE 1.037e-17
CC47765 ZN A1:2 2.702e-17
R14 M7:SRC M8:DRN 0.001 
CC47801 M7:SRC M7:GATE 4.59e-18
CC47756 M7:SRC A1:1 2.434e-17
CC47892 M7:SRC M8:GATE 3.088e-17
R15 M1:SRC M2:DRN 0.001 
CC47788 M1:SRC M2:GATE 5.1e-18
CC47816 M1:SRC A2:1 2.778e-17
CC47764 M1:SRC A1:2 2.407e-17
CC47902 M1:SRC M1:GATE 5.33e-18
C16 M5:SRC 0 4.48e-18
C17 ZN:1 0 1.3e-16
C18 M14:SRC 0 5.23e-18
C19 ZN:2 0 2.409e-17
C20 M3:SRC 0 4.47e-18
C21 M10:SRC 0 5.7e-18
C22 ZN 0 1.352e-17
C23 M7:SRC 0 5.29e-18
C24 M1:SRC 0 5.73e-18
R25 M15:GATE A1:1 111.3 
CC47839 M15:GATE M16:GATE 1.344e-17
CC47806 M15:GATE A2:1 7.33e-18
R26 M7:GATE A1:1 94.0755 
R27 A1 A1:1 35.4028 
R28 M6:GATE A1:1 180.614 
R29 A1:1 M14:GATE 213.685 
CC47897 A1:1 M8:GATE 5.66e-18
CC47843 A1:1 M16:GATE 1.022e-17
CC47836 A1:1 A2:2 9.97e-18
CC47820 A1:1 A2:1 2.28e-18
R30 A1 M14:GATE 477.612 
R31 M14:GATE M6:GATE 834.495 
CC47825 M14:GATE A2:2 4.1e-18
CC47808 M14:GATE A2:1 8.42e-18
CC47846 M14:GATE M13:GATE 1.325e-17
R32 M6:GATE A1 403.695 
CC47876 M6:GATE M5:GATE 2.69e-18
CC47829 M6:GATE A2:2 1.57e-18
R33 A1 A1:2 23.9592 
CC47880 A1 M5:GATE 4.97e-18
CC47888 A1 M4:GATE 8.85e-18
CC47834 A1 A2:2 1.42e-17
CC47818 A1 A2:1 7.074e-17
R34 M3:GATE A1:2 92.22 
R35 M2:GATE A1:2 145.96 
R36 M10:GATE A1:2 153.703 
R37 A1:2 M11:GATE 105.205 
CC47890 A1:2 M4:GATE 3.49e-18
CC47866 A1:2 M9:GATE 1.064e-17
CC47821 A1:2 A2:1 1.87e-18
CC47837 A1:2 A2:2 1.148e-17
CC47852 M11:GATE M12:GATE 1.335e-17
CC47809 M11:GATE A2:1 8.03e-18
R38 M10:GATE M2:GATE 650.036 
CC47899 M10:GATE M1:GATE 7.03e-18
CC47864 M10:GATE M9:GATE 1.299e-17
CC47811 M10:GATE A2:1 9.47e-18
CC47901 M2:GATE M1:GATE 2.37e-18
CC47886 M3:GATE M4:GATE 2.86e-18
CC47893 M7:GATE M8:GATE 2.49e-18
C39 M15:GATE 0 3.975e-17
C40 A1:1 0 1.247e-17
C41 M14:GATE 0 3.768e-17
C42 M6:GATE 0 3.626e-17
C43 A1 0 5.74e-18
C44 A1:2 0 1.152e-17
C45 M11:GATE 0 4.418e-17
C46 M10:GATE 0 3.831e-17
C47 M2:GATE 0 4.518e-17
C48 M3:GATE 0 3.988e-17
C49 M7:GATE 0 4.486e-17
R50 M1:GATE M9:GATE 511.536 
R51 M9:GATE A2:1 145.573 
R52 M1:GATE A2:1 131.279 
R53 A2 A2:1 0.50963 
R54 M8:GATE A2:1 132.458 
R55 A2:1 M16:GATE 142.679 
R56 M16:GATE M8:GATE 506.953 
R57 M13:GATE A2:2 104.675 
R58 M5:GATE A2:2 93.1916 
R59 A2 A2:2 22.1453 
R60 M4:GATE A2:2 142.907 
R61 A2:2 M12:GATE 148.548 
R62 M12:GATE M4:GATE 695.372 
C63 M9:GATE 0 9.263e-17
C64 A2:1 0 4.5293e-16
C65 M16:GATE 0 8.929e-17
C66 M8:GATE 0 3.472e-17
C67 M13:GATE 0 5.163e-17
C68 A2:2 0 2.006e-17
C69 M12:GATE 0 5.375e-17
C70 M4:GATE 0 3.347e-17
C71 A2 0 4.46e-18
C72 M1:GATE 0 5.624e-17
C73 M5:GATE 0 3.079e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
