.SUBCKT OAI21D1 A1 A2 B ZN
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.3e-07  SB=4.6e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M1:DRN vss nch L=6e-08 W=3.97e-07  AD=7.8e-14  AS=3.9e-14  PD=1.18e-06  PS=5.9e-07  SA=6.9e-07  SB=2e-07  NRD=1.346  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.6e-14  PD=5.9e-07  PS=1.12e-06  SA=1.7e-07  SB=7.2e-07  NRD=4.183  NRS=0.583  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE M4:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.5e-14  PD=7.2e-07  PS=7.3e-07  SA=4.3e-07  SB=4.6e-07  NRD=2.099  NRS=0.202  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 M5:DRN M5:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=1.04e-13  PD=7.2e-07  PS=1.44e-06  SA=6.9e-07  SB=2e-07  NRD=2.099  NRS=1.435  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M4:SRC M6:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.5e-14  AS=8.3e-14  PD=7.3e-07  PS=1.36e-06  SA=1.6e-07  SB=7.3e-07  NRD=0.202  NRS=0.532  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M1:DRN M3:SRC 60.7653 
CC92625 M1:DRN M5:GATE 1.34e-18
CC92662 M1:DRN ZN 7.787e-17
CC92633 M1:DRN A1 2.67e-17
CC92636 M1:DRN M1:GATE 1.06e-17
CC92670 M1:DRN M1:SRC 2.86e-18
CC92644 M1:DRN A2 5.76e-18
CC92628 M1:DRN M2:GATE 9.46e-18
CC92627 M1:DRN B 2.629e-17
CC92643 M3:SRC A2 5.504e-17
CC92668 M3:SRC M1:SRC 2.76e-18
CC92640 M3:SRC M6:GATE 1.83e-18
CC92647 M3:SRC M3:GATE 2.58e-18
C1 M1:DRN 0 1.174e-17
C2 M3:SRC 0 9.04e-17
R3 M4:GATE A1 151.386 
R4 A1 M1:GATE 117.651 
CC92631 A1 M5:GATE 1.394e-17
CC92646 A1 A2 2.311e-17
CC92634 A1 M2:GATE 5.68e-18
CC92635 A1 B 4.515e-17
CC92667 A1 ZN 3.906e-17
CC92641 A1 M6:GATE 2.46e-18
CC92656 A1 M5:DRN 2.05e-18
CC92676 A1 M4:SRC 1.07e-18
CC92674 A1 M1:SRC 2.475e-17
CC92650 A1 M3:GATE 3.99e-18
R5 M1:GATE M4:GATE 540.545 
CC92645 M1:GATE A2 1.31e-18
CC92637 M1:GATE M2:GATE 1.25e-18
CC92638 M1:GATE B 3.93e-18
CC92664 M1:GATE ZN 4.58e-18
CC92649 M1:GATE M3:GATE 6.78e-18
CC92671 M1:GATE M1:SRC 1.167e-17
CC92639 M4:GATE M6:GATE 1.327e-17
CC92642 M4:GATE A2 1.419e-17
CC92659 M4:GATE ZN 4.74e-18
CC92653 M4:GATE M5:DRN 2.831e-17
CC92629 M4:GATE M5:GATE 7.47e-18
CC92630 M4:GATE B 1.48e-18
C6 A1 0 7.03e-18
C7 M1:GATE 0 3.434e-17
C8 M4:GATE 0 4.707e-17
R9 M3:DRN M1:SRC 0.001 
R10 M1:SRC ZN 31.2654 
CC92673 M1:SRC A2 1.284e-17
CC92669 M1:SRC M3:GATE 1.68e-17
R11 ZN M5:DRN 30.9847 
CC92658 ZN M5:GATE 9.65e-18
CC92661 ZN M3:GATE 2.78e-18
CC92663 ZN M2:GATE 7.53e-18
CC92665 ZN B 7.998e-17
CC92666 ZN A2 6.29e-18
R12 M5:DRN M4:DRN 0.001 
CC92652 M5:DRN M5:GATE 2.869e-17
CC92655 M5:DRN B 6.53e-18
C13 M1:SRC 0 4.58e-18
C14 ZN 0 1.2943e-16
C15 M5:DRN 0 6.58e-18
R16 B M2:GATE 117.651 
R17 M2:GATE M5:GATE 540.545 
R18 M5:GATE B 151.386 
C19 M2:GATE 0 5.719e-17
C20 M5:GATE 0 7.388e-17
C21 B 0 2.54e-17
R22 M3:GATE A2 113.425 
R23 A2 M6:GATE 147.705 
R24 M6:GATE M3:GATE 500.395 
C25 A2 0 3.63e-17
C26 M6:GATE 0 1.0017e-16
C27 M3:GATE 0 3.383e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
