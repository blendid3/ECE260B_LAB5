.SUBCKT INVD16 I ZN
MMM20 M20:DRN M20:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.28e-06  SB=9.2e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 vdd M21:GATE M21:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.02e-06  SB=1.18e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.76e-06  SB=1.44e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 vdd M23:GATE M23:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.5e-06  SB=1.7e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 M24:DRN M24:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.24e-06  SB=1.96e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM25 vdd M25:GATE M25:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.98e-06  SB=2.22e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM26 M26:DRN M26:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.72e-06  SB=2.48e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM27 vdd M27:GATE M27:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.46e-06  SB=2.74e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM28 M28:DRN M28:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.2e-06  SB=3e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM29 vdd M29:GATE M29:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.4e-07  SB=3.26e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.72e-06  SB=2.48e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.46e-06  SB=2.74e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=4.04e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.2e-06  SB=3e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=3.78e-06  SB=4.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.4e-07  SB=3.26e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=3.54e-06  SB=6.6e-07  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=3.52e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.28e-06  SB=9.2e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vss M15:GATE M15:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=3.78e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.02e-06  SB=1.18e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.2e-14  PD=5.9e-07  PS=1.1e-06  SA=1.6e-07  SB=4.04e-06  NRD=4.141  NRS=0.462  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.76e-06  SB=1.44e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 vdd M17:GATE M17:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=4.04e-06  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.5e-06  SB=1.7e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M18:DRN M18:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=3.78e-06  SB=4.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.24e-06  SB=1.96e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vdd M19:GATE M19:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=3.54e-06  SB=6.6e-07  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.98e-06  SB=2.22e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM30 M30:DRN M30:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=3.52e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM31 vdd M31:GATE M31:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=3.78e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM32 M32:DRN M32:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=4.04e-06  NRD=2.057  NRS=0.427  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M25:SRC M26:DRN 0.001 
R1 M26:DRN ZN:1 14.9999 
CC9489 M26:DRN I:16 1.1e-17
CC9585 M26:DRN M25:GATE 4.499e-17
CC9582 M26:DRN M26:GATE 4.525e-17
R2 ZN ZN:1 0.104 
R3 M30:DRN ZN:1 53.4962 
R4 M18:DRN ZN:1 16.3621 
R5 M20:DRN ZN:1 16.1748 
R6 M22:DRN ZN:1 15.7153 
R7 M24:DRN ZN:1 14.9999 
R8 M28:DRN ZN:1 26.5881 
R9 ZN:1 ZN:2 0.64389 
CC9450 ZN:1 M20:GATE 1.05e-18
CC9458 ZN:1 M18:GATE 1.11e-18
CC9435 ZN:1 I:8 1.334e-17
CC9442 ZN:1 M22:GATE 1.14e-18
CC9399 ZN:1 I:1 1.206e-17
CC9411 ZN:1 I:4 1.5e-18
CC9415 ZN:1 I:5 5.76e-18
CC9544 ZN:1 M9:GATE 1.84e-18
CC9505 ZN:1 I:16 3.685e-17
CC9592 ZN:1 M24:GATE 4.55e-18
CC9588 ZN:1 M25:GATE 1.004e-17
CC9580 ZN:1 M27:GATE 1.53e-18
CC9596 ZN:1 M23:GATE 1.24e-18
R10 M32:DRN ZN:2 14.9999 
R11 M30:DRN ZN:2 21.0937 
R12 ZN:2 M28:DRN 35.664 
CC9445 ZN:2 M21:GATE 1.751e-17
CC9449 ZN:2 M20:GATE 1.749e-17
CC9453 ZN:2 M19:GATE 1.841e-17
CC9457 ZN:2 M18:GATE 1.701e-17
CC9460 ZN:2 M17:GATE 5.15e-18
CC9434 ZN:2 I:8 1.0025e-16
CC9441 ZN:2 M22:GATE 1.683e-17
CC9398 ZN:2 I:1 9.765e-17
CC9567 ZN:2 M30:GATE 1.855e-17
CC9563 ZN:2 M31:GATE 1.65e-17
CC9559 ZN:2 M32:GATE 5.11e-18
CC9504 ZN:2 I:16 4.194e-17
CC9595 ZN:2 M23:GATE 1.716e-17
CC9591 ZN:2 M24:GATE 1.535e-17
CC9587 ZN:2 M25:GATE 1.474e-17
CC9583 ZN:2 M26:GATE 1.679e-17
CC9579 ZN:2 M27:GATE 1.67e-17
CC9575 ZN:2 M28:GATE 1.853e-17
CC9571 ZN:2 M29:GATE 1.67e-17
CC9602 ZN:2 I 8.13e-18
R13 M28:DRN M27:SRC 0.001 
CC9427 M28:DRN I:8 1.58e-18
CC9488 M28:DRN I:16 1.114e-17
CC9577 M28:DRN M27:GATE 4.495e-17
CC9574 M28:DRN M28:GATE 4.554e-17
R14 M24:DRN M23:SRC 0.001 
CC9490 M24:DRN I:16 1.104e-17
CC9593 M24:DRN M23:GATE 4.485e-17
CC9590 M24:DRN M24:GATE 4.487e-17
R15 M21:SRC M22:DRN 0.001 
R16 M18:DRN M22:DRN 906.26 
R17 M22:DRN M20:DRN 1269.06 
CC9443 M22:DRN M21:GATE 4.484e-17
CC9390 M22:DRN I:1 1.57e-18
CC9440 M22:DRN M22:GATE 4.478e-17
CC9491 M22:DRN I:16 1.114e-17
R18 M19:SRC M20:DRN 0.001 
R19 M20:DRN M18:DRN 539.859 
CC9448 M20:DRN M20:GATE 4.454e-17
CC9451 M20:DRN M19:GATE 4.48e-17
CC9391 M20:DRN I:1 1.57e-18
CC9492 M20:DRN I:16 1.114e-17
R20 M18:DRN M17:SRC 0.001 
CC9456 M18:DRN M18:GATE 4.452e-17
CC9459 M18:DRN M17:GATE 4.586e-17
CC9392 M18:DRN I:1 1.5e-18
CC9493 M18:DRN I:16 1.098e-17
R21 M15:SRC M16:DRN 0.001 
R22 M14:DRN M16:DRN 524.507 
R23 M12:DRN M16:DRN 880.699 
R24 M16:DRN ZN:3 16.414 
CC9429 M16:DRN I:8 1.13e-18
CC9436 M16:DRN I:9 2.726e-17
CC9556 M16:DRN M15:GATE 4.59e-18
CC9494 M16:DRN I:16 1.614e-17
CC9516 M16:DRN M16:GATE 1.917e-17
CC9510 M16:DRN I:18 4.082e-17
R25 M8:DRN ZN:3 14.9999 
R26 M10:DRN ZN:3 14.9999 
R27 M14:DRN ZN:3 16.2126 
R28 M4:DRN ZN:3 16.2127 
R29 M6:DRN ZN:3 15.8221 
R30 ZN ZN:3 0.03813 
R31 M12:DRN ZN:3 15.8219 
R32 ZN:3 M2:DRN 16.4065 
CC9464 ZN:3 I:11 2.97e-18
CC9423 ZN:3 I:7 1.26e-18
CC9433 ZN:3 I:8 1.3056e-16
CC9397 ZN:3 I:1 1.3337e-16
CC9404 ZN:3 I:3 1.75e-18
CC9414 ZN:3 I:5 1.38e-18
CC9545 ZN:3 M10:GATE 1.56e-17
CC9543 ZN:3 M9:GATE 1.206e-17
CC9537 ZN:3 M13:GATE 1.406e-17
CC9534 ZN:3 M12:GATE 1.566e-17
CC9532 ZN:3 M1:GATE 3.98e-18
CC9529 ZN:3 M2:GATE 1.242e-17
CC9526 ZN:3 M3:GATE 1.469e-17
CC9523 ZN:3 M4:GATE 1.359e-17
CC9555 ZN:3 M15:GATE 1.376e-17
CC9552 ZN:3 M14:GATE 1.563e-17
CC9550 ZN:3 M11:GATE 1.444e-17
CC9483 ZN:3 I:15 3.12e-18
CC9478 ZN:3 I:14 2.84e-18
CC9473 ZN:3 I:13 2.5e-18
CC9520 ZN:3 M5:GATE 1.226e-17
CC9517 ZN:3 M6:GATE 1.345e-17
CC9515 ZN:3 M16:GATE 4.13e-18
CC9508 ZN:3 I:17 1.32e-18
CC9503 ZN:3 I:16 5.996e-17
CC9608 ZN:3 M7:GATE 4.72e-18
CC9606 ZN:3 M8:GATE 1.18e-17
CC9601 ZN:3 I 4.4e-18
R33 M4:DRN M2:DRN 524.271 
R34 M6:DRN M2:DRN 880.294 
R35 M2:DRN M1:SRC 0.001 
CC9396 M2:DRN I:1 1.08e-18
CC9400 M2:DRN I:2 4.129e-17
CC9533 M2:DRN M1:GATE 4.8e-18
CC9531 M2:DRN M2:GATE 4.59e-18
CC9482 M2:DRN I:15 4.014e-17
CC9501 M2:DRN I:16 1.614e-17
R36 M14:DRN M12:DRN 869.889 
R37 M12:DRN M11:SRC 0.001 
CC9422 M12:DRN I:7 3.848e-17
CC9431 M12:DRN I:8 1.37e-18
CC9416 M12:DRN I:6 3.795e-17
CC9536 M12:DRN M12:GATE 6.8e-18
CC9548 M12:DRN M11:GATE 7.29e-18
CC9496 M12:DRN I:16 1.643e-17
R38 M29:SRC M30:DRN 0.001 
CC9426 M30:DRN I:8 1.58e-18
CC9569 M30:DRN M29:GATE 4.495e-17
CC9566 M30:DRN M30:GATE 4.557e-17
CC9487 M30:DRN I:16 1.114e-17
R39 M31:SRC M32:DRN 0.001 
CC9425 M32:DRN I:8 1.55e-18
CC9560 M32:DRN M31:GATE 4.484e-17
CC9558 M32:DRN M32:GATE 4.595e-17
CC9486 M32:DRN I:16 1.105e-17
R40 M4:DRN M6:DRN 869.898 
R41 M6:DRN M5:SRC 0.001 
CC9462 M6:DRN I:11 4.077e-17
CC9394 M6:DRN I:1 1.07e-18
CC9403 M6:DRN I:3 3.756e-17
CC9522 M6:DRN M5:GATE 4.57e-18
CC9518 M6:DRN M6:GATE 7.52e-18
CC9499 M6:DRN I:16 1.677e-17
R42 M4:DRN M3:SRC 0.001 
CC9395 M4:DRN I:1 1.07e-18
CC9527 M4:DRN M3:GATE 4.57e-18
CC9524 M4:DRN M4:GATE 4.57e-18
CC9476 M4:DRN I:14 4.041e-17
CC9472 M4:DRN I:13 4.037e-17
CC9500 M4:DRN I:16 1.643e-17
R43 M14:DRN M13:SRC 0.001 
CC9467 M14:DRN I:12 4.067e-17
CC9430 M14:DRN I:8 1.37e-18
CC9538 M14:DRN M13:GATE 4.57e-18
CC9554 M14:DRN M14:GATE 4.57e-18
CC9507 M14:DRN I:17 4.077e-17
CC9495 M14:DRN I:16 1.643e-17
R44 M10:DRN M9:SRC 0.001 
CC9408 M10:DRN I:4 6.132e-17
CC9412 M10:DRN I:5 1.982e-17
CC9540 M10:DRN M9:GATE 5.98e-18
CC9547 M10:DRN M10:GATE 4.57e-18
CC9497 M10:DRN I:16 1.626e-17
R45 M8:DRN M7:SRC 0.001 
CC9413 M8:DRN I:5 4.075e-17
CC9498 M8:DRN I:16 5.008e-17
CC9611 M8:DRN M7:GATE 1.156e-17
CC9605 M8:DRN M8:GATE 4.57e-18
C46 M26:DRN 0 4.34e-18
C47 ZN:1 0 3.88e-18
C48 ZN:2 0 4.0406e-16
C49 M28:DRN 0 6.11e-18
C50 M24:DRN 0 4.34e-18
C51 M22:DRN 0 7.97e-18
C52 M20:DRN 0 1.569e-17
C53 M18:DRN 0 1.797e-17
C54 M16:DRN 0 7.38e-18
C55 ZN:3 0 3.9425e-16
C56 M2:DRN 0 7.26e-18
C57 M12:DRN 0 4.6e-18
C58 M30:DRN 0 6.63e-18
C59 M32:DRN 0 9.91e-18
C60 ZN 0 2.3e-19
C61 M6:DRN 0 4.66e-18
C62 M4:DRN 0 3.15e-18
C63 M14:DRN 0 4.64e-18
C64 M10:DRN 0 4.49e-18
C65 M8:DRN 0 4.49e-18
R66 M26:GATE I:4 111.3 
R67 M10:GATE I:4 94.0755 
R68 M25:GATE I:4 275.689 
R69 I:8 I:4 76.2668 
R70 I:6 I:4 30.4865 
R71 I:5 I:4 60.2341 
R72 I:4 M9:GATE 233.022 
R73 M25:GATE M9:GATE 1066.52 
R74 M9:GATE I:5 233.022 
R75 M8:GATE I:5 94.0755 
R76 M24:GATE I:5 111.3 
R77 M25:GATE I:5 275.689 
R78 I:5 I:16 24.3177 
R79 M23:GATE I:16 88.7752 
R80 M7:GATE I:16 94.0755 
R81 I:3 I:16 30.6013 
R82 I:16 I:1 65.6908 
R83 I:13 I:1 22 
R84 I:15 I:1 23.1442 
R85 I:2 I:1 23.385 
R86 I:14 I:1 22.6748 
R87 I:3 I:1 24.4481 
R88 I:1 I:11 17.8211 
R89 M21:GATE I:11 111.3 
R90 M5:GATE I:11 81.2035 
R91 I:13 I:11 22.4472 
R92 I:11 I:3 35.3042 
R93 M6:GATE I:3 94.0755 
R94 I:3 M22:GATE 111.3 
R95 M27:GATE I:6 111.3 
R96 M11:GATE I:6 94.0755 
R97 I:7 I:6 31.0275 
R98 I:6 I:8 24.2303 
R99 I:10 I:8 0.69247 
R100 I:7 I:8 29.3535 
R101 I:8 I:12 45.4767 
R102 I:10 I:12 29.8079 
R103 M13:GATE I:12 82.8124 
R104 M29:GATE I:12 100.037 
R105 I:17 I:12 21.9794 
R106 I:12 I:7 33.904 
R107 I:10 I:7 118.673 
R108 M28:GATE I:7 111.3 
R109 I:7 M12:GATE 94.0755 
R110 M30:GATE I:17 103.792 
R111 I:10 I:17 22 
R112 M14:GATE I:17 86.5669 
R113 I:17 I:18 21.5119 
R114 I:10 I:18 32.926 
R115 M15:GATE I:18 83.8364 
R116 M31:GATE I:18 101.061 
R117 I:9 I:18 22.3658 
R118 I:18 I 68.4613 
R119 I:10 I 0.70947 
R120 I I:9 34.0542 
R121 M16:GATE I:9 80.5597 
R122 I:10 I:9 64.0913 
R123 I:9 M32:GATE 97.7846 
R124 M3:GATE I:14 86.5669 
R125 I:13 I:14 21.0442 
R126 M19:GATE I:14 111.3 
R127 I:15 I:14 21.3057 
R128 I:14 I:2 2248.3 
R129 M1:GATE I:2 80.5597 
R130 I:15 I:2 22.0053 
R131 I:2 M17:GATE 111.3 
R132 M2:GATE I:15 83.8364 
R133 I:15 M18:GATE 111.3 
R134 M20:GATE I:13 111.3 
R135 I:13 M4:GATE 85.0652 
C136 M26:GATE 0 5.054e-17
C137 I:4 0 3.95e-18
C138 M9:GATE 0 3.261e-17
C139 I:5 0 1.04e-18
C140 I:16 0 1.437e-16
C141 I:1 0 3.426e-17
C142 I:11 0 7.35e-18
C143 I:3 0 4.02e-18
C144 M22:GATE 0 1.407e-17
C145 M27:GATE 0 3.512e-17
C146 I:6 0 3.36e-18
C147 I:8 0 1.42e-17
C148 I:12 0 4.59e-18
C149 I:7 0 2.8e-18
C150 M12:GATE 0 1.994e-17
C151 M25:GATE 0 4.482e-17
C152 M24:GATE 0 4.589e-17
C153 M30:GATE 0 4.109e-17
C154 I:17 0 4.49e-18
C155 I:18 0 3.61e-18
C156 I 0 6.754e-17
C157 I:9 0 3.337e-17
C158 M32:GATE 0 6.444e-17
C159 M29:GATE 0 3.465e-17
C160 M28:GATE 0 3.233e-17
C161 M8:GATE 0 3.179e-17
C162 M7:GATE 0 3.709e-17
C163 M23:GATE 0 4.801e-17
C164 M31:GATE 0 3.905e-17
C165 M13:GATE 0 2.296e-17
C166 M3:GATE 0 2.405e-17
C167 I:14 0 2.42e-18
C168 I:2 0 2.677e-17
C169 M17:GATE 0 7.14e-17
C170 M2:GATE 0 3.239e-17
C171 I:15 0 2.75e-18
C172 M18:GATE 0 2.468e-17
C173 M1:GATE 0 4.95e-17
C174 M14:GATE 0 2.854e-17
C175 M15:GATE 0 3.121e-17
C176 M10:GATE 0 3.448e-17
C177 M11:GATE 0 2.337e-17
C178 M19:GATE 0 1.809e-17
C179 I:13 0 2.83e-18
C180 M4:GATE 0 2.901e-17
C181 I:10 0 1.27e-17
C182 M5:GATE 0 2.237e-17
C183 M6:GATE 0 2.318e-17
C184 M16:GATE 0 2.793e-17
C185 M20:GATE 0 9.14e-18
C186 M21:GATE 0 1.508e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
