.SUBCKT OAI21D2 A1 A2 B ZN
MMM10 M9:SRC M10:GATE M10:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.6e-07  SB=9.4e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 M11:DRN M11:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=4e-07  SB=1.2e-06  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.567  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=8.3e-14  AS=4.7e-14  PD=1.36e-06  PS=7e-07  SA=1.6e-07  SB=1.44e-06  NRD=0.532  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.18e-06  SB=4.2e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M2:SRC M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.2e-07  SB=6.8e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE M4:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.6e-07  SB=9.4e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 M4:SRC M5:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=4e-07  SB=1.2e-06  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 vss M6:GATE M6:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=6.2e-14  PD=5.7e-07  PS=1.1e-06  SA=1.6e-07  SB=1.44e-06  NRD=7.648  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 M7:DRN M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.532  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M7:SRC M8:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.18e-06  SB=4.2e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.2e-07  SB=6.8e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M4:SRC M2:SRC 121.407 
R1 M6:SRC M2:SRC 124.303 
R2 M2:SRC M1:DRN 118.744 
CC92746 M2:SRC M6:GATE 2.23e-18
CC92740 M2:SRC M5:GATE 4.15e-18
CC92682 M2:SRC M4:GATE 4.68e-18
CC92683 M2:SRC M1:GATE 8.42e-18
CC92706 M2:SRC M1:SRC 5.48e-18
CC92704 M2:SRC M3:SRC 5.14e-18
CC92699 M2:SRC ZN 6.22e-18
CC92787 M2:SRC M3:GATE 3.5e-17
CC92777 M2:SRC M2:GATE 1.505e-17
CC92773 M2:SRC A2 1.02e-18
CC92752 M2:SRC A2:1 2.373e-17
R3 M4:SRC M1:DRN 124.417 
R4 M1:DRN M6:SRC 127.384 
CC92680 M1:DRN A1 2.483e-17
CC92684 M1:DRN M1:GATE 4.27e-18
CC92707 M1:DRN M1:SRC 1.01e-18
CC92701 M1:DRN ZN 1.3e-18
CC92716 M1:DRN B:1 6.17e-18
CC92772 M1:DRN A2 2.43e-18
R5 M6:SRC M4:SRC 118.639 
CC92733 M6:SRC B 1.07e-18
CC92713 M6:SRC B:1 2.862e-17
CC92696 M6:SRC ZN 8.767e-17
CC92678 M4:SRC A1 3.763e-17
CC92737 M4:SRC M5:GATE 9.18e-18
CC92681 M4:SRC M4:GATE 9.33e-18
CC92734 M4:SRC B 1.819e-17
CC92697 M4:SRC ZN 6.456e-17
CC92714 M4:SRC B:1 2.255e-17
CC92749 M4:SRC A2:1 4.57e-18
C6 M2:SRC 0 5.812e-17
C7 M1:DRN 0 9.59e-17
C8 M6:SRC 0 3.751e-17
C9 M4:SRC 0 9.88e-18
CC92709 M7:SRC A1 1.11e-18
CC92748 M9:SRC A2:1 1.08e-18
R10 A1 M4:GATE 121.354 
R11 M4:GATE M10:GATE 542.94 
CC92715 M4:GATE B:1 5.29e-18
CC92770 M4:GATE A2 3.81e-18
CC92738 M4:GATE M5:GATE 3.44e-18
CC92750 M4:GATE A2:1 7.68e-18
CC92784 M4:GATE M3:GATE 3.39e-18
CC92698 M4:GATE ZN 8.34e-18
R12 M10:GATE A1 147.094 
CC92712 M10:GATE B:1 1.082e-17
CC92758 M10:GATE M9:GATE 1.516e-17
CC92747 M10:GATE A2:1 5.55e-18
CC92726 M10:GATE M11:GATE 7.85e-18
CC92694 M10:GATE ZN 6.96e-18
CC92685 M10:GATE M10:SRC 3.04e-17
R13 M1:GATE A1 124.501 
R14 A1 M7:GATE 150.91 
CC92767 A1 M8:GATE 6.17e-18
CC92768 A1 A2 6.532e-17
CC92756 A1 A2:1 1.005e-17
CC92728 A1 M11:GATE 2.4e-18
CC92783 A1 M3:GATE 1.04e-18
CC92761 A1 M9:GATE 4.84e-18
CC92736 A1 B 3.03e-18
CC92693 A1 M7:DRN 1.74e-18
CC92687 A1 M10:SRC 5.89e-18
CC92708 A1 M1:SRC 3.72e-17
CC92702 A1 ZN 1.8202e-16
CC92705 A1 M3:SRC 3.052e-17
R15 M7:GATE M1:GATE 516.533 
CC92763 M7:GATE M8:GATE 1.429e-17
CC92695 M7:GATE ZN 7.54e-18
CC92690 M7:GATE M7:DRN 2.851e-17
CC92771 M1:GATE A2 1.25e-18
CC92779 M1:GATE M2:GATE 3.62e-18
CC92765 M1:GATE M8:GATE 5.72e-18
CC92754 M1:GATE A2:1 1.107e-17
CC92700 M1:GATE ZN 3.41e-18
C16 M4:GATE 0 2.891e-17
C17 M10:GATE 0 4.168e-17
C18 A1 0 1.498e-17
C19 M7:GATE 0 5.55e-17
C20 M1:GATE 0 3.303e-17
R21 M1:SRC M3:SRC 1027.49 
R22 M4:DRN M3:SRC 0.001 
R23 M3:SRC ZN 31.889 
CC92751 M3:SRC A2:1 3.763e-17
CC92774 M3:SRC A2 2.01e-18
CC92739 M3:SRC M5:GATE 1.63e-18
R24 M1:SRC ZN 32.8116 
R25 M10:SRC ZN 32.196 
R26 M12:DRN ZN 32.4196 
R27 ZN M7:DRN 33.6224 
CC92743 ZN M6:GATE 1.4e-18
CC92741 ZN M5:GATE 2.4e-18
CC92769 ZN A2 4.085e-17
CC92766 ZN M8:GATE 6.31e-18
CC92781 ZN M2:GATE 6.21e-18
CC92760 ZN M9:GATE 3.56e-18
CC92755 ZN A2:1 2.65e-18
CC92722 ZN M12:GATE 8.57e-18
CC92727 ZN M11:GATE 1.745e-17
CC92717 ZN B:1 9.79e-18
CC92735 ZN B 7.004e-17
R28 M10:SRC M7:DRN 1250.04 
R29 M7:DRN M12:DRN 1636.09 
R30 M12:DRN M10:SRC 1566.69 
CC92719 M12:DRN M12:GATE 2.83e-17
CC92729 M12:DRN B 1.87e-18
R31 M10:SRC M11:DRN 0.001 
CC92725 M10:SRC M11:GATE 2.833e-17
R32 M1:SRC M2:DRN 0.001 
CC92753 M1:SRC A2:1 4.35e-18
CC92778 M1:SRC M2:GATE 2.949e-17
C33 M3:SRC 0 1.9e-18
C34 ZN 0 1.4887e-16
C35 M7:DRN 0 3.096e-17
C36 M12:DRN 0 1.103e-17
C37 M10:SRC 0 9.74e-18
C38 M1:SRC 0 1.91e-18
R39 B:1 M5:GATE 130.664 
R40 M5:GATE M11:GATE 733.433 
R41 M11:GATE B:1 154.587 
R42 M6:GATE B:1 83.3024 
R43 M12:GATE B:1 111.3 
R44 B:1 B 22 
C45 M5:GATE 0 4.036e-17
C46 M11:GATE 0 4.825e-17
C47 B:1 0 2.942e-17
C48 B 0 1.351e-17
C49 M12:GATE 0 5.233e-17
C50 M6:GATE 0 4.383e-17
R51 M3:GATE A2:1 82.8124 
R52 M8:GATE A2:1 170.513 
R53 M2:GATE A2:1 144.124 
R54 M9:GATE A2:1 111.3 
R55 A2:1 A2 22.065 
R56 M2:GATE M8:GATE 591.409 
C57 M3:GATE 0 2.294e-17
C58 A2:1 0 3.592e-17
C59 M9:GATE 0 8.707e-17
C60 M2:GATE 0 1.577e-17
C61 M8:GATE 0 7.836e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
