.SUBCKT DFCSNQD4 D CP CDN SDN Q
MMM20 M19:SRC M20:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=5.1e-14  PD=5.9e-07  PS=7.99e-07  SA=3.08e-07  SB=2.005e-06  NRD=4.12  NRS=3.924  SCA=11.955  SCB=0.013  SCC=0.001 
MMM21 vss M21:GATE M12:SRC vss nch L=6e-08 W=2.17e-07  AD=2.8e-14  AS=2.1e-14  PD=4.31e-07  PS=4.1e-07  SA=4.45e-07  SB=2.29e-06  NRD=0.625  NRS=7.652  SCA=17.402  SCB=0.019  SCC=0.002 
MMM22 vdd M22:GATE M22:SRC vdd pch L=6e-08 W=3.54e-07  AD=4.5e-14  AS=3.5e-14  PD=9.6e-07  PS=5.5e-07  SA=1.35e-07  SB=2.55e-06  NRD=1.551  NRS=3.039  SCA=12.653  SCB=0.014  SCC=0.001 
MMM23 M22:SRC M23:GATE vdd vdd pch L=6e-08 W=3.55e-07  AD=3.5e-14  AS=4.3e-14  PD=5.5e-07  PS=5.99e-07  SA=3.96e-07  SB=2.29e-06  NRD=3.039  NRS=0.603  SCA=12.653  SCB=0.014  SCC=0.001 
MMM24 M24:DRN M24:GATE vdd vdd pch L=6e-08 W=1.55e-07  AD=2.6e-14  AS=2e-14  PD=6.5e-07  PS=4.15e-07  SA=1.75e-07  SB=6.2e-07  NRD=1.195  NRS=0.955  SCA=14.652  SCB=0.018  SCC=0.001 
MMM25 M25:DRN M25:GATE M25:SRC vdd pch L=6e-08 W=1.87e-07  AD=2.9e-14  AS=2.1e-14  PD=6.22e-07  PS=3.71e-07  SA=5.9e-07  SB=1.8e-07  NRD=0.9  NRS=0.667  SCA=6.102  SCB=0.006  SCC=0.0001158 
MMM26 M26:DRN M26:GATE M26:SRC vdd pch L=6e-08 W=1.53e-07  AD=2.6e-14  AS=1.7e-14  PD=6.5e-07  PS=3.35e-07  SA=4.25e-07  SB=1.75e-07  NRD=1.195  NRS=0.755  SCA=20.527  SCB=0.023  SCC=0.003 
MMM27 M27:DRN M27:GATE M26:SRC vdd pch L=6e-08 W=2.8e-07  AD=4.4e-14  AS=3.1e-14  PD=8.9e-07  PS=6.25e-07  SA=1.55e-07  SB=2.28e-07  NRD=0.66  NRS=14.264  SCA=14.603  SCB=0.016  SCC=0.002 
MMM28 vdd M28:GATE M28:SRC vdd pch L=6e-08 W=4.82e-07  AD=6.7e-14  AS=4.8e-14  PD=1.36e-06  PS=6.8e-07  SA=4.96e-07  SB=1.34e-07  NRD=0.524  NRS=2.258  SCA=10.228  SCB=0.011  SCC=0.0008915 
MMM29 M28:SRC M29:GATE vdd vdd pch L=6e-08 W=4.84e-07  AD=4.8e-14  AS=6.4e-14  PD=6.8e-07  PS=1.329e-06  SA=2e-07  SB=3.97e-07  NRD=2.258  NRS=0.731  SCA=7.816  SCB=0.008  SCC=0.0004769 
MMM40 M39:SRC M40:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.7e-14  PD=7.2e-07  PS=7.4e-07  SA=9.91e-07  SB=1.465e-06  NRD=2.099  NRS=0.689  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM41 vdd M41:GATE M41:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.7e-14  AS=5.2e-14  PD=7.4e-07  PS=7.2e-07  SA=6.83e-07  SB=1.745e-06  NRD=0.689  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM42 M41:SRC M42:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.4e-14  PD=7.2e-07  PS=8.91e-07  SA=3.57e-07  SB=2.005e-06  NRD=2.099  NRS=1.145  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.4e-14  AS=3.5e-14  PD=1.11e-06  PS=5.7e-07  SA=4e-07  SB=1.65e-07  NRD=0.575  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=6.2e-14  PD=5.7e-07  PS=1.1e-06  SA=1.6e-07  SB=4.05e-07  NRD=7.648  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=2.12e-07  AD=1.5e-14  AS=2.3e-14  PD=3.5e-07  PS=4.39e-07  SA=8.38e-07  SB=4.34e-07  NRD=24.729  NRS=0.538  SCA=12.705  SCB=0.015  SCC=0.001 
MMM12 M12:DRN M12:GATE M12:SRC vss nch L=6e-08 W=2.1e-07  AD=3.9e-14  AS=2.1e-14  PD=7.9e-07  PS=4.1e-07  SA=1.85e-07  SB=2.55e-06  NRD=0.935  NRS=7.652  SCA=17.402  SCB=0.019  SCC=0.002 
MMM2 M1:DRN M2:GATE vss vss nch L=6e-08 W=2.18e-07  AD=1.5e-14  AS=2.9e-14  PD=3.5e-07  PS=5.37e-07  SA=5.23e-07  SB=6.79e-07  NRD=24.729  NRS=0.881  SCA=14.662  SCB=0.017  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.97e-07  AD=6.6e-14  AS=3.9e-14  PD=1.12e-06  PS=5.9e-07  SA=2.276e-06  SB=1.7e-07  NRD=1.416  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=1.5e-07  AD=1.3e-14  AS=1.3e-14  PD=3.2e-07  PS=3.2e-07  SA=6.85e-07  SB=1.356e-06  NRD=22.667  NRS=22.667  SCA=20.648  SCB=0.023  SCC=0.003 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.011e-06  SB=4.3e-07  NRD=4.183  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE M4:SRC vss nch L=6e-08 W=3.94e-07  AD=3.8e-14  AS=4.4e-14  PD=6.62e-07  PS=8.52e-07  SA=2.67e-07  SB=2.17e-07  NRD=8.254  NRS=10.891  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vss M15:GATE M15:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.746e-06  SB=6.9e-07  NRD=4.537  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 M1:SRC M5:GATE M5:SRC vss nch L=6.1e-08 W=2.32e-07  AD=2.5e-14  AS=2.5e-14  PD=4.81e-07  PS=5.21e-07  SA=5.54e-07  SB=2.7e-07  NRD=5.114  NRS=11.621  SCA=16.515  SCB=0.019  SCC=0.002 
MMM16 M16:DRN M16:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.8e-14  PD=5.9e-07  PS=5.85e-07  SA=1.478e-06  SB=9.5e-07  NRD=4.183  NRS=5.314  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 vss M6:GATE M4:DRN vss nch L=6e-08 W=3.1e-07  AD=5e-14  AS=3e-14  PD=9.4e-07  PS=5.18e-07  SA=1.65e-07  SB=3.78e-07  NRD=0.65  NRS=1.015  SCA=7.268  SCB=0.008  SCC=0.0002566 
MMM17 vss M17:GATE M17:SRC vss nch L=6e-08 W=3.96e-07  AD=3.8e-14  AS=3.9e-14  PD=5.85e-07  PS=5.9e-07  SA=1.213e-06  SB=1.205e-06  NRD=5.314  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vss M7:GATE M3:DRN vss nch L=6e-08 W=1.59e-07  AD=2.1e-14  AS=1.3e-14  PD=3.83e-07  PS=3.2e-07  SA=9.2e-07  SB=1.124e-06  NRD=1.048  NRS=22.667  SCA=20.648  SCB=0.023  SCC=0.003 
MMM18 M17:SRC M18:GATE M18:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4.3e-14  PD=5.9e-07  PS=6.1e-07  SA=9.37e-07  SB=1.465e-06  NRD=4.12  NRS=1.112  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M8:DRN M8:GATE M5:SRC vss nch L=6e-08 W=1.55e-07  AD=2.6e-14  AS=1.7e-14  PD=6.5e-07  PS=3.39e-07  SA=9.56e-07  SB=1.75e-07  NRD=1.195  NRS=0.746  SCA=20.622  SCB=0.023  SCC=0.003 
MMM19 M18:SRC M19:GATE M19:SRC vss nch L=6e-08 W=3.9e-07  AD=4.3e-14  AS=3.9e-14  PD=6.1e-07  PS=5.9e-07  SA=6.28e-07  SB=1.745e-06  NRD=1.112  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 M4:SRC M9:GATE M3:SRC vss nch L=6e-08 W=1.56e-07  AD=1.7e-14  AS=1.3e-14  PD=3.28e-07  PS=3.2e-07  SA=4.48e-07  SB=1.588e-06  NRD=0.762  NRS=22.667  SCA=20.648  SCB=0.023  SCC=0.003 
MMM30 M25:DRN M30:GATE vdd vdd pch L=6e-08 W=1.58e-07  AD=2.4e-14  AS=2e-14  PD=5.18e-07  PS=4.15e-07  SA=1.3e-07  SB=2.5e-07  NRD=1.072  NRS=0.955  SCA=3.346  SCB=0.002  SCC=4.515e-06 
MMM31 M25:SRC M31:GATE M31:SRC vdd pch L=6e-08 W=4.95e-07  AD=5.9e-14  AS=3.5e-14  PD=1.019e-06  PS=6.35e-07  SA=3.3e-07  SB=1.91e-07  NRD=10.371  NRS=14.773  SCA=8.408  SCB=0.009  SCC=0.0005868 
MMM32 M31:SRC M32:GATE vdd vdd pch L=6e-08 W=4.99e-07  AD=3.5e-14  AS=6.4e-14  PD=6.35e-07  PS=1.25e-06  SA=1.3e-07  SB=4.12e-07  NRD=14.773  NRS=1.814  SCA=8.408  SCB=0.009  SCC=0.0005868 
MMM33 M33:DRN M33:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=8.1e-14  AS=4.7e-14  PD=1.36e-06  PS=7e-07  SA=4e-07  SB=1.57e-07  NRD=0.53  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM34 vdd M34:GATE M34:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=8.3e-14  PD=7e-07  PS=1.36e-06  SA=1.6e-07  SB=3.97e-07  NRD=6.61  NRS=0.532  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM35 vdd M35:GATE M35:SRC vdd pch L=6e-08 W=5.24e-07  AD=8.8e-14  AS=5.2e-14  PD=1.38e-06  PS=7.2e-07  SA=2.323e-06  SB=1.7e-07  NRD=0.44  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM36 M36:DRN M36:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.06e-06  SB=4.3e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM37 vdd M37:GATE M37:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.795e-06  SB=6.9e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM38 M38:DRN M38:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.1e-14  PD=7.2e-07  PS=7.15e-07  SA=1.529e-06  SB=9.5e-07  NRD=2.099  NRS=3.552  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM39 vdd M39:GATE M39:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.1e-14  AS=5.2e-14  PD=7.15e-07  PS=7.2e-07  SA=1.265e-06  SB=1.205e-06  NRD=3.552  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 Q M35:SRC 30.3359 
R1 M35:SRC M36:DRN 0.001 
CC67505 M35:SRC M36:GATE 2.782e-17
CC67484 M35:SRC N_12:2 1.108e-17
CC67507 M35:SRC M35:GATE 2.829e-17
R2 Q M37:SRC 30.4618 
R3 M37:SRC M38:DRN 0.001 
CC67466 M37:SRC N_12:1 1.53e-18
CC67497 M37:SRC M38:GATE 2.834e-17
CC67501 M37:SRC M37:GATE 2.768e-17
CC67483 M37:SRC N_12:2 1.109e-17
R4 M15:SRC Q 30.3174 
R5 Q M13:SRC 30.2242 
CC67555 Q M16:GATE 3.08e-18
CC67559 Q M18:SRC 1.41e-18
CC67550 Q M15:GATE 1.115e-17
CC67546 Q M14:GATE 9.43e-18
CC67544 Q M13:GATE 8.61e-18
CC67488 Q N_12:2 4.433e-17
CC67494 Q N_12:3 4.03e-18
CC67503 Q M37:GATE 1.716e-17
CC67498 Q M38:GATE 4.56e-18
CC67506 Q M36:GATE 1.248e-17
CC67509 Q M35:GATE 7.58e-18
CC67477 Q N_12:1 9.004e-17
R6 M13:SRC M14:DRN 0.001 
CC67545 M13:SRC M13:GATE 8.53e-18
CC67487 M13:SRC N_12:2 1.44e-17
CC67493 M13:SRC N_12:3 4.772e-17
CC67508 M13:SRC M35:GATE 2.66e-18
R7 M15:SRC M16:DRN 0.001 
CC67554 M15:SRC M16:GATE 5.3e-18
CC67548 M15:SRC M15:GATE 2.67e-18
CC67492 M15:SRC N_12:3 1.285e-17
CC67486 M15:SRC N_12:2 5.245e-17
CC67474 M15:SRC N_12:1 1.33e-18
C8 M35:SRC 0 6.78e-18
C9 M37:SRC 0 5.3e-18
C10 Q 0 1.4532e-16
C11 M13:SRC 0 5.74e-18
C12 M15:SRC 0 5.74e-18
CC67580 M3:SRC N_19:1 1.41e-18
CC67258 M4:DRN D 1.6e-18
CC67386 M17:SRC CDN:1 1.17e-18
CC67394 M12:SRC CDN:2 1.49e-18
R13 M22:GATE M12:GATE 357.824 
R14 M12:GATE SDN 99.9317 
CC67266 M12:GATE N_26:1 7.27e-18
CC67530 M12:GATE M23:GATE 1.41e-18
CC67248 M12:GATE M12:DRN 1.631e-17
CC67538 M12:GATE M21:GATE 9.28e-18
CC67247 M12:GATE M26:DRN 4.04e-18
R15 SDN M22:GATE 130.423 
CC67274 SDN N_26:1 1.25e-18
CC67282 SDN M26:GATE 1.56e-18
CC67244 SDN M22:SRC 9.399e-17
CC67243 SDN M26:DRN 2.14e-18
CC67532 SDN M23:GATE 9.52e-18
CC67245 SDN M12:DRN 2.314e-17
R16 M22:GATE M28:GATE 536.624 
CC67470 M22:GATE N_12:1 4.95e-18
CC67529 M22:GATE M23:GATE 4e-18
CC67242 M22:GATE M22:SRC 2.395e-17
CC67241 M22:GATE M26:DRN 1.299e-17
R17 M28:GATE M1:GATE 182.85 
CC67617 M28:GATE M28:SRC 3.151e-17
CC67276 M28:GATE M26:GATE 1.25e-18
CC67254 M28:GATE M4:SRC 4.89e-18
CC67589 M28:GATE M27:DRN 3.55e-18
CC67251 M28:GATE M26:DRN 1.55e-18
CC67250 M28:GATE M29:GATE 8.12e-18
CC67288 M28:GATE M5:GATE 3.94e-18
CC67632 M28:GATE M1:SRC 9.46e-18
CC67567 M28:GATE N_19:1 5.02e-18
CC67467 M28:GATE N_12:1 3.9e-18
CC67273 M1:GATE N_26:1 9.75e-18
CC67594 M1:GATE M27:DRN 2.07e-18
CC67257 M1:GATE M2:GATE 2.582e-17
CC67638 M1:GATE M1:SRC 2.209e-17
CC67582 M1:GATE N_19:1 8.17e-18
C18 M12:GATE 0 1.646e-17
C19 SDN 0 2.14e-17
C20 M22:GATE 0 9.382e-17
C21 M28:GATE 0 2.2297e-16
C22 M1:GATE 0 1.555e-17
R23 M22:SRC M26:DRN 118.59 
R24 M12:DRN M26:DRN 122.992 
R25 M26:DRN M8:DRN 122.51 
CC67289 M26:DRN M5:GATE 1.11e-18
CC67441 M26:DRN M26:SRC 1.88e-18
CC67427 M26:DRN N_30:2 5.62e-18
CC67390 M26:DRN CDN 3.44e-18
CC67391 M26:DRN CDN:2 3.83e-18
CC67334 M26:DRN M8:GATE 2.8e-18
CC67277 M26:DRN M26:GATE 3.647e-17
CC67264 M26:DRN N_26:1 5.592e-17
R26 M22:SRC M8:DRN 125.058 
R27 M8:DRN M12:DRN 117.933 
CC67442 M8:DRN M26:SRC 1.14e-18
CC67432 M8:DRN N_30:2 9.484e-17
CC67280 M8:DRN M26:GATE 5.34e-18
CC67292 M8:DRN M5:GATE 1.71e-18
CC67397 M8:DRN CDN:2 1.96e-18
CC67336 M8:DRN M8:GATE 3.191e-17
CC67269 M8:DRN N_26:1 2.718e-17
R28 M12:DRN M22:SRC 125.55 
CC67430 M12:DRN N_30:2 5.643e-17
CC67387 M12:DRN CDN:1 7.21e-18
CC67290 M12:DRN M5:GATE 2.48e-18
CC67395 M12:DRN CDN:2 5.37e-18
CC67267 M12:DRN N_26:1 1.37e-17
CC67475 M12:DRN N_12:1 3.51e-18
CC67428 M22:SRC N_30:2 1.563e-17
CC67528 M22:SRC M23:GATE 1.129e-17
CC67469 M22:SRC N_12:1 2.148e-17
C29 M26:DRN 0 2.223e-17
C30 M8:DRN 0 4.99e-18
C31 M12:DRN 0 3.863e-17
C32 M22:SRC 0 2.75e-18
R33 M25:SRC M4:SRC 76.4371 
R34 M2:GATE M4:SRC 232.391 
R35 M4:SRC M29:GATE 417.899 
CC67296 M4:SRC M9:GATE 1.64e-18
CC67366 M4:SRC M25:GATE 7.26e-18
CC67328 M4:SRC N_28:2 1.55e-18
CC67405 M4:SRC M7:GATE 1.733e-17
CC67403 M4:SRC M24:GATE 5.75e-18
CC67268 M4:SRC N_26:1 8.43e-18
CC67270 M4:SRC N_26:1 5.06e-18
CC67619 M4:SRC M28:SRC 1.4e-17
CC67239 M4:SRC D 9.495e-17
CC67294 M4:SRC M9:GATE 3.89e-17
CC67633 M4:SRC M1:SRC 1e-18
CC67237 M4:SRC M31:GATE 9.51e-18
CC67234 M4:SRC M24:DRN 1.965e-17
CC67233 M4:SRC M25:DRN 1.912e-17
CC67628 M4:SRC M3:GATE 1.372e-17
R36 M25:SRC M29:GATE 432.97 
R37 M29:GATE M2:GATE 319.562 
CC67322 M29:GATE N_28:2 2.22e-18
CC67350 M29:GATE N_28:1 4.38e-18
CC67400 M29:GATE M24:GATE 7.01e-18
CC67262 M29:GATE N_26:1 3.609e-17
CC67566 M29:GATE N_19:1 8.51e-18
CC67616 M29:GATE M28:SRC 2.106e-17
CC67605 M29:GATE M30:GATE 1.1e-18
R38 M2:GATE M25:SRC 240.775 
CC67398 M2:GATE CDN:2 1.07e-18
CC67272 M2:GATE N_26:1 2e-18
CC67581 M2:GATE N_19:1 6.274e-17
CC67320 M25:SRC N_28:2 2.702e-17
CC67348 M25:SRC N_28:1 1.74e-18
CC67363 M25:SRC M25:GATE 1.463e-17
CC67306 M25:SRC N_28:1 3.14e-17
CC67240 M25:SRC M4:GATE 1.94e-18
CC67564 M25:SRC N_19:1 5.949e-17
CC67238 M25:SRC D 4.08e-18
CC67261 M25:SRC N_26:1 9.907e-17
CC67235 M25:SRC M31:GATE 2.79e-17
C39 M4:SRC 0 1.243e-17
C40 M29:GATE 0 4.504e-17
C41 M2:GATE 0 2.292e-17
C42 M25:SRC 0 8.1e-18
R43 M24:DRN M25:DRN 60.6736 
CC67402 M24:DRN M24:GATE 3.179e-17
CC67310 M24:DRN N_28:1 1.21e-18
CC67610 M24:DRN M30:GATE 3.416e-17
CC67365 M24:DRN M25:GATE 1.75e-18
CC67572 M24:DRN N_19:1 5.748e-17
CC67326 M24:DRN N_28:2 3.34e-18
CC67404 M24:DRN M7:GATE 1.37e-18
CC67325 M25:DRN N_28:2 2.43e-18
CC67570 M25:DRN N_19:1 1.32e-18
CC67364 M25:DRN M25:GATE 3.415e-17
CC67608 M25:DRN M30:GATE 2.305e-17
CC67626 M25:DRN M3:GATE 4.51e-18
CC67309 M25:DRN N_28:1 6.117e-17
CC67351 M25:DRN N_28:1 3.43e-18
CC67401 M25:DRN M24:GATE 3.56e-18
CC67321 M25:DRN N_28:2 2.48e-18
C44 M24:DRN 0 1.192e-17
C45 M25:DRN 0 1.542e-17
R46 M4:GATE D 124.105 
R47 D M31:GATE 142.349 
CC67275 D N_26:1 6.535e-17
CC67299 D M9:GATE 3.32e-18
CC67285 D M32:GATE 5.5e-18
CC67383 D M6:GATE 1.301e-17
CC67314 D N_28:1 1.839e-17
R48 M31:GATE M4:GATE 531.699 
CC67283 M31:GATE M32:GATE 2.12e-17
CC67362 M31:GATE M25:GATE 3.79e-18
CC67347 M31:GATE N_28:1 3.08e-18
CC67319 M31:GATE N_28:2 3.15e-18
CC67305 M31:GATE N_28:1 2e-18
CC67381 M4:GATE M6:GATE 4.26e-18
CC67297 M4:GATE M9:GATE 2.12e-18
CC67271 M4:GATE N_26:1 2.391e-17
C49 D 0 1.257e-17
C50 M31:GATE 0 3.798e-17
C51 M4:GATE 0 3.113e-17
R52 M11:GATE CP 120.685 
R53 CP M34:GATE 146.49 
CC67374 CP M10:GATE 1.833e-17
CC67369 CP M11:SRC 3.625e-17
CC67355 CP N_28:1 2.344e-17
CC67359 CP M34:SRC 6.15e-18
CC67315 CP N_28:1 6.286e-17
R54 M34:GATE M11:GATE 536.415 
CC67302 M34:GATE N_28:1 9.48e-18
CC67357 M34:GATE M34:SRC 2.803e-17
CC67339 M34:GATE M33:GATE 1.457e-17
CC67344 M34:GATE N_28:1 7.7e-18
CC67371 M11:GATE M10:GATE 9.98e-18
CC67311 M11:GATE N_28:1 9.36e-18
CC67360 M11:GATE M34:SRC 1.5e-18
C55 CP 0 1.165e-17
C56 M34:GATE 0 5.269e-17
C57 M11:GATE 0 4.255e-17
R58 N_26:1 M26:GATE 254.457 
R59 M26:GATE M5:GATE 3651.45 
CC67426 M26:GATE N_30:2 8.49e-18
CC67440 M26:GATE M26:SRC 3.305e-17
CC67330 M26:GATE M27:GATE 2.01e-18
CC67333 M26:GATE M8:GATE 5.96e-18
R60 M9:GATE M5:GATE 4534.85 
R61 M5:GATE N_26:1 77.9633 
CC67433 M5:GATE N_30:2 5.18e-18
CC67337 M5:GATE M8:GATE 3.19e-18
CC67593 M5:GATE M27:DRN 2.08e-18
CC67458 M5:GATE M5:SRC 3.553e-17
CC67332 M5:GATE M27:GATE 2.53e-18
CC67579 M5:GATE N_19:1 5.07e-18
CC67636 M5:GATE M1:SRC 2.076e-17
R62 M32:GATE N_26:1 178.048 
R63 M10:DRN N_26:1 15.0688 
R64 M9:GATE N_26:1 87.6391 
R65 N_26:1 M33:DRN 30.6592 
CC67639 N_26:1 M1:SRC 1.034e-17
CC67435 N_26:1 N_30:2 2.373e-17
CC67343 N_26:1 M33:GATE 1.328e-17
CC67338 N_26:1 M8:GATE 5.89e-18
CC67459 N_26:1 M5:SRC 1.24e-18
CC67585 N_26:1 N_19:1 3.644e-17
CC67316 N_26:1 N_28:1 1.2161e-16
CC67630 N_26:1 M3:GATE 5.62e-18
CC67384 N_26:1 M6:GATE 1.508e-17
CC67375 N_26:1 M10:GATE 5.67e-18
CC67356 N_26:1 N_28:1 2.28e-18
CC67303 M33:DRN N_28:1 3.371e-17
CC67345 M33:DRN N_28:1 1.97e-18
CC67627 M9:GATE M3:GATE 8.03e-18
CC67573 M9:GATE N_19:1 8.18e-18
CC67312 M10:DRN N_28:1 8.48e-18
CC67378 M10:DRN M6:GATE 4.66e-18
CC67372 M10:DRN M10:GATE 5.886e-17
CC67304 M32:GATE N_28:1 5.19e-18
CC67346 M32:GATE N_28:1 4.27e-18
C66 M26:GATE 0 1.446e-17
C67 M5:GATE 0 3.117e-17
C68 N_26:1 0 3.671e-16
C69 M33:DRN 0 2.612e-17
C70 M9:GATE 0 2.602e-17
C71 M10:DRN 0 2.697e-17
C72 M32:GATE 0 3.267e-17
R73 M10:GATE M33:GATE 538.382 
R74 M33:GATE N_28:1 149.446 
R75 N_28:2 N_28:1 1.31542 
R76 M34:SRC N_28:1 30.1961 
R77 M10:GATE N_28:1 126.551 
R78 N_28:1 M11:SRC 31.9919 
CC67584 N_28:1 N_19:1 1.213e-17
CC67613 N_28:1 M30:GATE 1.36e-18
CC67621 N_28:1 M28:SRC 1.42e-18
CC67612 N_28:1 M30:GATE 5.5e-18
R79 M11:SRC M10:GATE 5104.04 
R80 M10:GATE M6:GATE 253.87 
R81 N_28:2 M27:GATE 81.0663 
R82 M27:GATE M8:GATE 134.941 
CC67590 M27:GATE M27:DRN 1.288e-17
CC67568 M27:GATE N_19:1 2.11e-18
CC67425 M27:GATE N_30:2 3.12e-18
CC67454 M27:GATE M5:SRC 1.096e-17
CC67439 M27:GATE M26:SRC 2.118e-17
CC67431 M8:GATE N_30:2 8.14e-18
CC67456 M8:GATE M5:SRC 2.353e-17
R83 N_28:2 M25:GATE 72.1458 
CC67586 N_28:2 N_19:1 7.998e-17
CC67615 N_28:2 M30:GATE 5.46e-18
CC67596 N_28:2 M27:DRN 2.913e-17
CC67444 N_28:2 M26:SRC 1.236e-17
CC67436 N_28:2 N_30:2 2.702e-17
CC67624 N_28:2 M28:SRC 7.98e-18
CC67607 M25:GATE M30:GATE 2.48e-18
C84 M33:GATE 0 1.971e-17
C85 N_28:1 0 2.6463e-16
C86 M11:SRC 0 1.958e-17
C87 M10:GATE 0 7.254e-17
C88 M6:GATE 0 7.676e-17
C89 M27:GATE 0 2.675e-17
C90 M8:GATE 0 7.26e-18
C91 M34:SRC 0 1.308e-17
C92 N_28:2 0 1.2988e-16
C93 M25:GATE 0 1.309e-17
R94 M42:GATE CDN:1 149.276 
R95 M20:GATE CDN:1 123.572 
R96 M17:GATE CDN:1 119.675 
R97 M39:GATE CDN:1 153.991 
R98 CDN:1 CDN 0.23833 
CC67481 CDN:1 N_12:1 7.862e-17
CC67423 CDN:1 M40:GATE 4.2e-18
CC67417 CDN:1 M41:GATE 6.95e-18
CC67411 CDN:1 N_30:1 2.886e-17
CC67453 CDN:1 M19:GATE 3.85e-18
CC67449 CDN:1 M18:GATE 1.124e-17
CC67438 CDN:1 N_30:2 5.607e-17
CC67561 CDN:1 M18:SRC 9.77e-18
CC67542 CDN:1 M21:GATE 1.042e-17
CC67535 CDN:1 M23:GATE 1.06e-17
CC67523 CDN:1 M39:SRC 1.041e-17
CC67516 CDN:1 M41:SRC 2.005e-17
CC67499 CDN:1 M38:GATE 1.8e-18
CC67489 CDN:1 N_12:2 1.937e-17
CC67434 CDN N_30:2 4.013e-17
CC67414 CDN M41:GATE 3.77e-18
CC67410 CDN N_30:1 2.69e-18
CC67514 CDN M41:SRC 2.6e-18
R99 M20:GATE CDN:2 691.648 
R100 CDN:2 M7:GATE 109.975 
CC67461 CDN:2 M5:SRC 2.33e-18
CC67452 CDN:2 M19:GATE 6.76e-18
CC67641 CDN:2 M1:SRC 2.78e-18
CC67541 CDN:2 M21:GATE 3.16e-18
R101 M7:GATE M24:GATE 129.849 
CC67629 M7:GATE M3:GATE 5.57e-18
CC67578 M7:GATE N_19:1 7.79e-18
CC67609 M24:GATE M30:GATE 2.27e-18
CC67571 M24:GATE N_19:1 1.869e-17
R102 M39:GATE M17:GATE 522.779 
CC67419 M39:GATE M40:GATE 6.5e-18
CC67408 M39:GATE N_30:1 2.34e-18
CC67465 M39:GATE N_12:1 2.115e-17
CC67520 M39:GATE M39:SRC 2.94e-17
CC67496 M39:GATE M38:GATE 1.381e-17
CC67485 M17:GATE N_12:2 1.33e-17
CC67447 M17:GATE M18:GATE 4.28e-18
CC67473 M17:GATE N_12:1 9.54e-18
CC67521 M17:GATE M39:SRC 3.07e-18
CC67553 M17:GATE M16:GATE 3.34e-18
R103 M20:GATE M42:GATE 554.351 
CC67409 M20:GATE N_30:1 9.78e-18
CC67450 M20:GATE M19:GATE 2.98e-18
CC67424 M42:GATE N_30:2 5.67e-18
CC67407 M42:GATE N_30:1 4.55e-18
CC67462 M42:GATE N_12:1 6.46e-18
CC67525 M42:GATE M23:GATE 1.33e-18
CC67510 M42:GATE M41:SRC 9.68e-18
C104 CDN:1 0 7.42e-17
C105 CDN:2 0 3.7665e-16
C106 M7:GATE 0 4.578e-17
C107 M24:GATE 0 2.588e-17
C108 M39:GATE 0 3.383e-17
C109 M17:GATE 0 2.141e-17
C110 M20:GATE 0 8.055e-17
C111 M42:GATE 0 3.226e-17
R112 M41:GATE N_30:1 104.675 
CC67511 M41:GATE M41:SRC 2.917e-17
CC67463 M41:GATE N_12:1 7.03e-18
R113 M19:GATE N_30:1 100.7 
R114 N_30:2 N_30:1 51.2697 
R115 M18:GATE N_30:1 239.445 
R116 N_30:1 M40:GATE 248.895 
CC67562 N_30:1 M18:SRC 4.236e-17
CC67517 N_30:1 M41:SRC 1.07e-18
CC67490 N_30:1 N_12:2 3.31e-18
R117 N_30:2 M40:GATE 328.721 
R118 M40:GATE M18:GATE 786.841 
CC67556 M40:GATE M18:SRC 2.6e-18
CC67464 M40:GATE N_12:1 6.79e-18
CC67519 M40:GATE M39:SRC 2.947e-17
R119 M18:GATE N_30:2 316.237 
CC67558 M18:GATE M18:SRC 7.58e-18
CC67472 M18:GATE N_12:1 5.91e-18
R120 M5:SRC N_30:2 30.9024 
R121 N_30:2 M26:SRC 29.9999 
CC67515 N_30:2 M41:SRC 6.23e-18
CC67560 N_30:2 M18:SRC 9.02e-18
CC67534 N_30:2 M23:GATE 5.35e-18
CC67631 N_30:2 M3:GATE 4.75e-18
CC67598 N_30:2 M27:DRN 2.93e-18
CC67588 N_30:2 N_19:1 5.834e-17
CC67522 N_30:2 M39:SRC 1.51e-18
CC67480 N_30:2 N_12:1 1.3945e-16
CC67592 M5:SRC M27:DRN 1.19e-18
CC67575 M5:SRC N_19:1 1.85e-18
CC67471 M19:GATE N_12:1 3.77e-18
C122 M41:GATE 0 2.677e-17
C123 N_30:1 0 2.291e-17
C124 M40:GATE 0 3.501e-17
C125 M18:GATE 0 3.196e-17
C126 N_30:2 0 7.239e-17
C127 M26:SRC 0 1.106e-17
C128 M5:SRC 0 5.49e-18
C129 M19:GATE 0 2.685e-17
R130 M39:SRC N_12:2 1240.34 
R131 M38:GATE N_12:2 111.3 
R132 M16:GATE N_12:2 82.3623 
R133 N_12:1 N_12:2 25.2424 
R134 M18:SRC N_12:2 479.522 
R135 N_12:3 N_12:2 64.6546 
R136 M15:GATE N_12:2 250.123 
R137 N_12:2 M37:GATE 295.921 
R138 N_12:3 M37:GATE 263.489 
R139 M37:GATE M15:GATE 1019.34 
R140 M15:GATE N_12:3 222.713 
R141 M36:GATE N_12:3 111.3 
R142 M14:GATE N_12:3 94.0755 
R143 M35:GATE N_12:3 164.389 
R144 N_12:3 M13:GATE 138.947 
R145 M13:GATE M35:GATE 635.948 
R146 M39:SRC M18:SRC 1752.77 
R147 M18:SRC N_12:1 35.6708 
R148 M39:SRC N_12:1 31.9293 
R149 M41:SRC N_12:1 29.9999 
R150 N_12:1 M23:GATE 98.6676 
R151 M23:GATE M21:GATE 159 
C152 N_12:2 0 3.455e-17
C153 M37:GATE 0 5.967e-17
C154 M15:GATE 0 3.121e-17
C155 N_12:3 0 1.369e-17
C156 M13:GATE 0 2.574e-17
C157 M35:GATE 0 7.868e-17
C158 M18:SRC 0 1.932e-17
C159 N_12:1 0 2.3744e-16
C160 M23:GATE 0 2.14e-17
C161 M21:GATE 0 4.031e-17
C162 M14:GATE 0 2.773e-17
C163 M16:GATE 0 2.256e-17
C164 M38:GATE 0 2.375e-17
C165 M41:SRC 0 6.45e-18
C166 M36:GATE 0 6.164e-17
C167 M39:SRC 0 6.43e-18
R168 N_19:1 M30:GATE 230.835 
R169 M30:GATE M3:GATE 528.598 
R170 M3:GATE N_19:1 86.6249 
R171 M28:SRC N_19:1 30.5038 
R172 M27:DRN N_19:1 30.3335 
R173 N_19:1 M1:SRC 30.4926 
C174 M30:GATE 0 3.649e-17
C175 M3:GATE 0 4.22e-18
C176 N_19:1 0 2.94e-17
C177 M1:SRC 0 2.8e-18
C178 M27:DRN 0 9.13e-18
C179 M28:SRC 0 4.47e-18
.ENDS
*.SCALE METER 
.GLOBAL VSS VDD
