.SUBCKT MUX2D0 I0 I1 S Z
MMM10 M8:SRC M10:GATE M9:DRN vdd pch L=6e-08 W=2.6e-07  AD=1.9e-14  AS=2.6e-14  PD=4.05e-07  PS=4.6e-07  SA=6e-07  SB=6.05e-07  NRD=26.117  NRS=4.054  SCA=7.615  SCB=0.009  SCC=0.0002993 
MMM11 M9:SRC M11:GATE vdd vdd pch L=6e-08 W=2.66e-07  AD=2.8e-14  AS=5.1e-14  PD=5.25e-07  PS=7.49e-07  SA=2.29e-07  SB=4.01e-07  NRD=0.41  NRS=0.911  SCA=12.084  SCB=0.014  SCC=0.001 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=2.02e-07  AD=3.4e-14  AS=1.8e-14  PD=7.4e-07  PS=3.75e-07  SA=6.8e-07  SB=1.75e-07  NRD=0.947  NRS=14.653  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=2.56e-07  AD=4.1e-14  AS=4.9e-14  PD=8.3e-07  PS=7.21e-07  SA=1.65e-07  SB=2.31e-07  NRD=0.741  NRS=0.93  SCA=4.146  SCB=0.003  SCC=2.287e-05 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=2.02e-07  AD=1.8e-14  AS=1.4e-14  PD=3.75e-07  PS=3.35e-07  SA=4.33e-07  SB=4.15e-07  NRD=14.653  NRS=26.632  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM3 M2:SRC M3:GATE M3:SRC vss nch L=6e-08 W=2.02e-07  AD=1.4e-14  AS=4e-14  PD=3.35e-07  PS=6.35e-07  SA=2.25e-07  SB=6.15e-07  NRD=26.632  NRS=1.045  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=1.95e-07  AD=3.5e-14  AS=2e-14  PD=7.5e-07  PS=3.95e-07  SA=1.8e-07  SB=7.55e-07  NRD=0.972  NRS=8.262  SCA=15.959  SCB=0.019  SCC=0.002 
MMM5 M3:SRC M5:GATE M5:SRC vss nch L=6e-08 W=2.02e-07  AD=4e-14  AS=1.9e-14  PD=6.35e-07  PS=3.9e-07  SA=6.95e-07  SB=2.25e-07  NRD=1.045  NRS=9.773  SCA=15.959  SCB=0.019  SCC=0.002 
MMM6 M5:SRC M6:GATE vss vss nch L=6e-08 W=1.95e-07  AD=1.9e-14  AS=2e-14  PD=3.9e-07  PS=3.95e-07  SA=4.4e-07  SB=4.89e-07  NRD=9.773  NRS=8.262  SCA=15.959  SCB=0.019  SCC=0.002 
MMM7 M7:DRN M7:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=4.2e-14  AS=2.3e-14  PD=8.4e-07  PS=4.4e-07  SA=1.072e-06  SB=1.6e-07  NRD=0.704  NRS=12.397  SCA=7.615  SCB=0.009  SCC=0.0002993 
MMM8 vdd M8:GATE M8:SRC vdd pch L=6e-08 W=2.65e-07  AD=2.3e-14  AS=1.9e-14  PD=4.4e-07  PS=4.05e-07  SA=8.21e-07  SB=4e-07  NRD=12.397  NRS=26.117  SCA=7.615  SCB=0.009  SCC=0.0002993 
MMM9 M9:DRN M9:GATE M9:SRC vdd pch L=6e-08 W=2.62e-07  AD=2.6e-14  AS=2.8e-14  PD=4.6e-07  PS=5.25e-07  SA=2.87e-07  SB=8.65e-07  NRD=4.054  NRS=0.41  SCA=7.615  SCB=0.009  SCC=0.0002993 
R0 M7:DRN Z 30.4298 
CC2801 M7:DRN M9:DRN 2.799e-17
CC2797 M7:DRN M7:GATE 8.49e-18
R1 Z M1:DRN 30.4396 
CC2829 Z M2:GATE 1.6e-18
CC2822 Z I1 2.41e-17
CC2807 Z M3:SRC 4.595e-17
CC2804 Z M1:GATE 4.65e-18
CC2799 Z M7:GATE 1.802e-17
CC2805 M1:DRN M1:GATE 2.406e-17
CC2798 M1:DRN M7:GATE 7.19e-18
C2 M7:DRN 0 2.06e-17
C3 Z 0 6.557e-17
C4 M1:DRN 0 1.791e-17
CC2882 M5:SRC M4:GATE 1.39e-18
CC2796 M5:SRC I0 1.62e-18
R5 M9:DRN M3:SRC 51.3585 
R6 M3:SRC M7:GATE 141.419 
CC2851 M3:SRC M5:GATE 1.636e-17
CC2843 M3:SRC M12:DRN 2.022e-17
CC2834 M3:SRC M10:GATE 1.433e-17
CC2893 M3:SRC M3:GATE 1.394e-17
CC2894 M3:SRC M3:GATE 2.082e-17
CC2886 M3:SRC M4:GATE 1.535e-17
CC2820 M3:SRC I1 5.359e-17
CC2844 M3:SRC M12:DRN 9.37e-18
CC2852 M3:SRC M5:GATE 1.656e-17
CC2810 M3:SRC I0 1.88e-17
CC2809 M3:SRC M6:GATE 1.72e-18
CC2819 M3:SRC I1 5.26e-18
R7 M9:DRN M7:GATE 270.779 
R8 M7:GATE M1:GATE 224.454 
CC2842 M7:GATE M12:DRN 2.614e-17
CC2824 M7:GATE M2:GATE 2.17e-18
CC2817 M7:GATE I1 1.812e-17
CC2827 M1:GATE M2:GATE 3.04e-18
CC2814 M1:GATE M8:GATE 1.719e-17
CC2875 M9:DRN S 1.19e-18
CC2866 M9:DRN M9:GATE 3.513e-17
CC2847 M9:DRN M5:GATE 2.451e-17
CC2840 M9:DRN M12:DRN 1.172e-17
CC2832 M9:DRN M10:GATE 3.96e-17
CC2823 M9:DRN M2:GATE 1.07e-18
CC2889 M9:DRN M3:GATE 1.179e-17
CC2811 M9:DRN M8:GATE 1.943e-17
CC2800 M9:DRN M11:GATE 3.49e-18
CC2802 M9:DRN M6:GATE 1.34e-18
C9 M3:SRC 0 9.92e-17
C10 M7:GATE 0 6.989e-17
C11 M1:GATE 0 2.749e-17
C12 M9:DRN 0 1.48e-17
R13 M2:GATE M8:GATE 653.046 
R14 M8:GATE I1 133.459 
CC2848 M8:GATE M5:GATE 1.644e-17
CC2841 M8:GATE M12:DRN 8.16e-18
R15 I1 M2:GATE 155.242 
CC2897 I1 M3:GATE 7.8e-18
CC2853 I1 M5:GATE 1.028e-17
CC2836 I1 M10:GATE 4.5e-18
CC2895 M2:GATE M3:GATE 1.177e-17
CC2887 M2:GATE M4:GATE 1.14e-18
C16 M8:GATE 0 2.53e-17
C17 I1 0 2.574e-17
C18 M2:GATE 0 3.545e-17
R19 M4:DRN M12:DRN 72.3596 
R20 M12:DRN M10:GATE 194.331 
CC2846 M12:DRN I0 2.856e-17
CC2838 M12:DRN M11:GATE 5.71e-18
CC2879 M12:DRN M4:GATE 1.706e-17
CC2856 M12:DRN M12:GATE 3.397e-17
CC2873 M12:DRN S 1.59e-18
CC2863 M12:DRN M9:GATE 1.82e-17
R21 M5:GATE M10:GATE 252.281 
R22 M10:GATE M4:DRN 199.512 
CC2837 M10:GATE I0 9.65e-18
CC2890 M10:GATE M3:GATE 3.48e-18
CC2867 M10:GATE M9:GATE 6.48e-18
CC2877 M4:DRN S 7.307e-17
CC2885 M4:DRN M4:GATE 2.458e-17
CC2850 M5:GATE M6:GATE 9.71e-18
CC2883 M5:GATE M4:GATE 3.51e-18
C23 M12:DRN 0 5.532e-17
C24 M10:GATE 0 9.664e-17
C25 M4:DRN 0 1.3579e-16
C26 M5:GATE 0 4.38e-18
CC2858 M9:SRC M12:GATE 1.13e-18
CC2865 M9:SRC M9:GATE 2.02e-18
CC2794 M9:SRC M11:GATE 1.58e-18
R27 M6:GATE M11:GATE 331.902 
R28 M11:GATE I0 112.207 
CC2874 M11:GATE S 1.342e-17
CC2857 M11:GATE M12:GATE 2.18e-18
CC2864 M11:GATE M9:GATE 1.276e-17
R29 I0 M6:GATE 108.676 
CC2888 I0 M4:GATE 6.15e-18
CC2878 I0 S 4.445e-17
CC2872 I0 M9:GATE 1.92e-18
CC2862 I0 M12:GATE 1.85e-18
CC2881 M6:GATE M4:GATE 6.35e-18
C30 M11:GATE 0 3.284e-17
C31 I0 0 4.636e-17
C32 M6:GATE 0 4.351e-17
R33 M3:GATE M4:GATE 389.814 
R34 M12:GATE M4:GATE 564.979 
R35 M4:GATE S 101.767 
R36 S M12:GATE 184.85 
R37 M12:GATE M9:GATE 324.625 
C38 M3:GATE 0 5.778e-17
C39 M4:GATE 0 1.3459e-16
C40 S 0 5.809e-17
C41 M12:GATE 0 1.25e-16
C42 M9:GATE 0 3.16e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
