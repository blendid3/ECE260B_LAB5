.SUBCKT DFCSNQD2 D CP CDN SDN Q
MMM20 vdd M20:GATE M20:SRC vdd pch L=6e-08 W=3.54e-07  AD=4.5e-14  AS=3.5e-14  PD=9.6e-07  PS=5.5e-07  SA=1.35e-07  SB=1.96e-06  NRD=1.551  NRS=3.039  SCA=12.653  SCB=0.014  SCC=0.001 
MMM21 M20:SRC M21:GATE vdd vdd pch L=6e-08 W=3.55e-07  AD=3.5e-14  AS=4.1e-14  PD=5.5e-07  PS=5.91e-07  SA=3.96e-07  SB=1.7e-06  NRD=3.039  NRS=0.598  SCA=12.653  SCB=0.014  SCC=0.001 
MMM22 M22:DRN M22:GATE M22:SRC vdd pch L=6e-08 W=1.87e-07  AD=2.9e-14  AS=2.1e-14  PD=6.22e-07  PS=3.71e-07  SA=5.9e-07  SB=1.8e-07  NRD=0.9  NRS=0.667  SCA=6.102  SCB=0.006  SCC=0.0001158 
MMM23 M23:DRN M23:GATE vdd vdd pch L=6e-08 W=1.55e-07  AD=2.6e-14  AS=2e-14  PD=6.5e-07  PS=4.15e-07  SA=1.75e-07  SB=6.2e-07  NRD=1.195  NRS=0.955  SCA=14.652  SCB=0.018  SCC=0.001 
MMM24 M24:DRN M24:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=4.1e-14  AS=2.3e-14  PD=8.4e-07  PS=4.4e-07  SA=4e-07  SB=1.58e-07  NRD=0.698  NRS=12.397  SCA=5.267  SCB=0.005  SCC=7.585e-05 
MMM25 M25:DRN M25:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=4.2e-14  AS=2.3e-14  PD=8.4e-07  PS=4.4e-07  SA=1.6e-07  SB=3.98e-07  NRD=0.704  NRS=12.397  SCA=5.267  SCB=0.005  SCC=7.585e-05 
MMM26 M26:DRN M26:GATE M26:SRC vdd pch L=6e-08 W=1.53e-07  AD=2.6e-14  AS=1.7e-14  PD=6.5e-07  PS=3.35e-07  SA=4.25e-07  SB=1.75e-07  NRD=1.195  NRS=0.755  SCA=20.527  SCB=0.023  SCC=0.003 
MMM27 M27:DRN M27:GATE M26:SRC vdd pch L=6e-08 W=2.8e-07  AD=4.4e-14  AS=3.1e-14  PD=8.9e-07  PS=6.25e-07  SA=1.55e-07  SB=2.28e-07  NRD=0.66  NRS=14.264  SCA=14.603  SCB=0.016  SCC=0.002 
MMM28 vdd M28:GATE M28:SRC vdd pch L=6e-08 W=4.84e-07  AD=6.4e-14  AS=4.8e-14  PD=1.329e-06  PS=6.8e-07  SA=2e-07  SB=3.97e-07  NRD=0.731  NRS=2.258  SCA=7.816  SCB=0.008  SCC=0.0004769 
MMM29 M22:DRN M29:GATE vdd vdd pch L=6e-08 W=1.58e-07  AD=2.4e-14  AS=2e-14  PD=5.18e-07  PS=4.15e-07  SA=1.3e-07  SB=2.5e-07  NRD=1.072  NRS=0.955  SCA=3.346  SCB=0.002  SCC=4.515e-06 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=2.04e-07  AD=3.4e-14  AS=1.8e-14  PD=7.4e-07  PS=3.75e-07  SA=4.15e-07  SB=1.75e-07  NRD=0.947  NRS=14.653  SCA=8.121  SCB=0.009  SCC=0.0003028 
MMM11 M11:DRN M11:GATE vss vss nch L=6e-08 W=2.04e-07  AD=3.4e-14  AS=1.8e-14  PD=7.4e-07  PS=3.75e-07  SA=1.75e-07  SB=4.15e-07  NRD=0.947  NRS=14.653  SCA=8.121  SCB=0.009  SCC=0.0003028 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=2.18e-07  AD=1.5e-14  AS=2.9e-14  PD=3.5e-07  PS=5.37e-07  SA=5.23e-07  SB=6.79e-07  NRD=24.729  NRS=0.881  SCA=14.662  SCB=0.017  SCC=0.001 
MMM12 M12:DRN M12:GATE M12:SRC vss nch L=6e-08 W=2.1e-07  AD=3.9e-14  AS=2.1e-14  PD=7.9e-07  PS=4.1e-07  SA=1.85e-07  SB=1.96e-06  NRD=0.935  NRS=7.652  SCA=17.402  SCB=0.019  SCC=0.002 
MMM2 M2:DRN M2:GATE M2:SRC vss nch L=6e-08 W=1.5e-07  AD=1.3e-14  AS=1.3e-14  PD=3.2e-07  PS=3.2e-07  SA=6.85e-07  SB=1.356e-06  NRD=22.667  NRS=22.667  SCA=20.648  SCB=0.023  SCC=0.003 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.97e-07  AD=5.1e-14  AS=3.9e-14  PD=1.04e-06  PS=5.9e-07  SA=1.715e-06  SB=1.3e-07  NRD=1.615  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=3.94e-07  AD=4.4e-14  AS=3.8e-14  PD=8.52e-07  PS=6.62e-07  SA=2.71e-07  SB=2.17e-07  NRD=10.891  NRS=8.254  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.7e-14  PD=5.9e-07  PS=5.8e-07  SA=1.447e-06  SB=3.9e-07  NRD=4.141  NRS=6.091  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M3:DRN M4:GATE M2:DRN vss nch L=6e-08 W=1.56e-07  AD=1.7e-14  AS=1.3e-14  PD=3.28e-07  PS=3.2e-07  SA=4.48e-07  SB=1.588e-06  NRD=0.762  NRS=22.667  SCA=20.648  SCB=0.023  SCC=0.003 
MMM15 vss M15:GATE M15:SRC vss nch L=6e-08 W=3.97e-07  AD=3.7e-14  AS=3.9e-14  PD=5.8e-07  PS=5.9e-07  SA=1.187e-06  SB=6.4e-07  NRD=6.091  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 M1:DRN M5:GATE M5:SRC vss nch L=6e-08 W=2.12e-07  AD=1.5e-14  AS=2.3e-14  PD=3.5e-07  PS=4.39e-07  SA=8.38e-07  SB=4.34e-07  NRD=24.729  NRS=0.538  SCA=12.705  SCB=0.015  SCC=0.001 
MMM16 M15:SRC M16:GATE M16:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4e-14  PD=5.9e-07  PS=5.95e-07  SA=9.1e-07  SB=9e-07  NRD=4.12  NRS=3.415  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 vss M6:GATE M3:SRC vss nch L=6e-08 W=3.1e-07  AD=5.3e-14  AS=3e-14  PD=9.6e-07  PS=5.18e-07  SA=1.75e-07  SB=3.78e-07  NRD=0.676  NRS=1.015  SCA=7.268  SCB=0.008  SCC=0.0002566 
MMM17 M16:SRC M17:GATE M17:SRC vss nch L=6e-08 W=3.9e-07  AD=4e-14  AS=3.9e-14  PD=5.95e-07  PS=5.9e-07  SA=6.16e-07  SB=1.165e-06  NRD=3.415  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 M5:SRC M7:GATE M7:SRC vss nch L=6.1e-08 W=2.32e-07  AD=2.5e-14  AS=2.5e-14  PD=4.81e-07  PS=5.21e-07  SA=5.54e-07  SB=2.7e-07  NRD=5.114  NRS=11.621  SCA=16.515  SCB=0.019  SCC=0.002 
MMM18 M17:SRC M18:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4.9e-14  PD=5.9e-07  PS=7.86e-07  SA=2.94e-07  SB=1.425e-06  NRD=4.12  NRS=5.497  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 vss M8:GATE M2:SRC vss nch L=6e-08 W=1.59e-07  AD=2.1e-14  AS=1.3e-14  PD=3.83e-07  PS=3.2e-07  SA=9.2e-07  SB=1.124e-06  NRD=1.048  NRS=22.667  SCA=20.648  SCB=0.023  SCC=0.003 
MMM19 vss M19:GATE M12:SRC vss nch L=6e-08 W=2.17e-07  AD=2.6e-14  AS=2.1e-14  PD=4.24e-07  PS=4.1e-07  SA=4.45e-07  SB=1.7e-06  NRD=0.608  NRS=7.652  SCA=17.402  SCB=0.019  SCC=0.002 
MMM9 M9:DRN M9:GATE M7:SRC vss nch L=6e-08 W=1.55e-07  AD=2.6e-14  AS=1.7e-14  PD=6.5e-07  PS=3.39e-07  SA=9.56e-07  SB=1.75e-07  NRD=1.195  NRS=0.746  SCA=20.622  SCB=0.023  SCC=0.003 
MMM30 M22:SRC M30:GATE M30:SRC vdd pch L=6e-08 W=4.95e-07  AD=5.9e-14  AS=3.5e-14  PD=1.019e-06  PS=6.35e-07  SA=3.3e-07  SB=1.91e-07  NRD=10.371  NRS=14.773  SCA=8.408  SCB=0.009  SCC=0.0005868 
MMM31 M28:SRC M31:GATE vdd vdd pch L=6e-08 W=4.82e-07  AD=4.8e-14  AS=6.7e-14  PD=6.8e-07  PS=1.36e-06  SA=4.96e-07  SB=1.34e-07  NRD=2.258  NRS=0.524  SCA=10.228  SCB=0.011  SCC=0.0008915 
MMM32 M30:SRC M32:GATE vdd vdd pch L=6e-08 W=4.99e-07  AD=3.5e-14  AS=6.4e-14  PD=6.35e-07  PS=1.25e-06  SA=1.3e-07  SB=4.12e-07  NRD=14.773  NRS=1.814  SCA=8.408  SCB=0.009  SCC=0.0005868 
MMM33 vdd M33:GATE M33:SRC vdd pch L=6e-08 W=5.24e-07  AD=6.8e-14  AS=5.2e-14  PD=1.3e-06  PS=7.2e-07  SA=1.765e-06  SB=1.3e-07  NRD=1.865  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM34 M34:DRN M34:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.9e-14  PD=7.2e-07  PS=7.1e-07  SA=1.498e-06  SB=3.9e-07  NRD=2.057  NRS=4.571  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM35 vdd M35:GATE M35:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.9e-14  AS=5.2e-14  PD=7.1e-07  PS=7.2e-07  SA=1.239e-06  SB=6.4e-07  NRD=4.571  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM36 M35:SRC M36:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.3e-14  PD=7.2e-07  PS=7.25e-07  SA=9.64e-07  SB=9e-07  NRD=2.099  NRS=1.517  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM37 vdd M37:GATE M37:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.3e-14  AS=5.2e-14  PD=7.25e-07  PS=7.2e-07  SA=6.71e-07  SB=1.165e-06  NRD=1.517  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM38 M37:SRC M38:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.1e-14  PD=7.2e-07  PS=8.79e-07  SA=3.43e-07  SB=1.425e-06  NRD=2.099  NRS=3.178  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M13:SRC M14:DRN 0.001 
R1 M14:DRN Q 15.2603 
CC67046 M14:DRN M13:GATE 2.018e-17
CC67052 M14:DRN M14:GATE 1.737e-17
CC66997 M14:DRN N_15:2 7.266e-17
CC66986 M14:DRN N_15:1 1.97e-18
R2 Q M34:DRN 15.3786 
CC67056 Q M16:SRC 2.23e-18
CC67049 Q M14:GATE 4.49e-18
CC67047 Q M13:GATE 1.532e-17
CC67008 Q M33:GATE 2.729e-17
CC67004 Q M34:GATE 5.41e-18
CC66998 Q N_15:2 1.592e-17
CC66989 Q N_15:1 1.0183e-16
R3 M34:DRN M33:SRC 0.001 
CC66995 M34:DRN N_15:2 1.408e-17
CC67007 M34:DRN M33:GATE 5.024e-17
CC67003 M34:DRN M34:GATE 4.922e-17
CC66977 M34:DRN N_15:1 2.42e-18
C4 M14:DRN 0 1.016e-17
C5 Q 0 8.382e-17
C6 M34:DRN 0 1.301e-17
CC67077 M2:DRN N_8:1 1.41e-18
CC66760 M3:SRC D 1.6e-18
CC66889 M3:SRC M6:GATE 3.25e-18
CC66897 M15:SRC CDN:1 1.16e-18
CC66905 M12:SRC CDN:2 1.48e-18
R7 SDN M20:GATE 130.423 
R8 M12:GATE M20:GATE 357.824 
R9 M20:GATE M31:GATE 536.624 
CC67029 M20:GATE M21:GATE 4e-18
CC66744 M20:GATE M26:DRN 1.294e-17
CC66745 M20:GATE M20:SRC 2.453e-17
CC66981 M20:GATE N_15:1 3.32e-18
R10 M31:GATE M5:GATE 182.85 
CC66788 M31:GATE M7:GATE 3.94e-18
CC66777 M31:GATE M26:GATE 1.27e-18
CC67129 M31:GATE M5:SRC 9.46e-18
CC67113 M31:GATE M28:SRC 3.147e-17
CC66754 M31:GATE M26:DRN 1.55e-18
CC66753 M31:GATE M28:GATE 8.12e-18
CC66978 M31:GATE N_15:1 5.99e-18
CC67060 M31:GATE N_8:1 4.96e-18
CC67085 M31:GATE M27:DRN 3.54e-18
CC66770 M5:GATE N_40:1 8.88e-18
CC67090 M5:GATE M27:DRN 2.05e-18
CC67133 M5:GATE M5:SRC 2.21e-17
CC66759 M5:GATE M1:GATE 2.733e-17
CC66758 M5:GATE M3:DRN 3.5e-18
CC67074 M5:GATE N_8:1 7.85e-18
R11 M12:GATE SDN 99.9317 
CC66767 M12:GATE N_40:1 2.95e-18
CC67039 M12:GATE M19:GATE 9.3e-18
CC67030 M12:GATE M21:GATE 1.71e-18
CC66751 M12:GATE M12:DRN 1.937e-17
CC66750 M12:GATE M26:DRN 4.19e-18
CC66782 SDN M26:GATE 5.82e-18
CC66775 SDN N_40:1 1.25e-18
CC67032 SDN M21:GATE 9.25e-18
CC66748 SDN M12:DRN 1.995e-17
CC66747 SDN M20:SRC 9.391e-17
CC66746 SDN M26:DRN 2.07e-18
C12 M20:GATE 0 9.524e-17
C13 M31:GATE 0 2.2631e-16
C14 M5:GATE 0 1.091e-17
C15 M12:GATE 0 1.659e-17
C16 SDN 0 2.012e-17
R17 M20:SRC M12:DRN 125.549 
R18 M26:DRN M12:DRN 122.992 
R19 M12:DRN M9:DRN 117.932 
CC66941 M12:DRN N_44:2 7.763e-17
CC66791 M12:DRN M7:GATE 2.48e-18
CC66768 M12:DRN N_40:1 1.374e-17
CC66987 M12:DRN N_15:1 3.56e-18
CC66898 M12:DRN CDN:1 7.22e-18
CC66906 M12:DRN CDN:2 5.37e-18
R20 M20:SRC M9:DRN 125.059 
R21 M9:DRN M26:DRN 122.51 
CC66943 M9:DRN N_44:2 6.747e-17
CC66792 M9:DRN M7:GATE 1.32e-18
CC66953 M9:DRN M26:SRC 1.14e-18
CC66769 M9:DRN N_40:1 5.688e-17
CC66907 M9:DRN CDN:2 1.96e-18
CC66837 M9:DRN M9:GATE 3.197e-17
CC66781 M9:DRN M26:GATE 5.34e-18
R22 M26:DRN M20:SRC 118.59 
CC66835 M26:DRN M9:GATE 2.86e-18
CC66902 M26:DRN CDN:2 3.88e-18
CC66952 M26:DRN M26:SRC 1.49e-18
CC66795 M26:DRN M4:GATE 1.11e-18
CC66938 M26:DRN N_44:2 1.054e-17
CC66789 M26:DRN M7:GATE 2.063e-17
CC66766 M26:DRN N_40:1 1.172e-17
CC66778 M26:DRN M26:GATE 3.052e-17
CC66901 M26:DRN CDN 3.48e-18
CC66939 M20:SRC N_44:2 1.678e-17
CC67028 M20:SRC M21:GATE 1.129e-17
CC66980 M20:SRC N_15:1 2.148e-17
C23 M12:DRN 0 1.452e-17
C24 M9:DRN 0 2.85e-18
C25 M26:DRN 0 4.596e-17
C26 M20:SRC 0 1.2e-18
R27 M11:GATE M25:GATE 639.968 
R28 M25:GATE CP 162.973 
CC66809 M25:GATE N_42:1 1.181e-17
CC66846 M25:GATE N_42:1 8.49e-18
CC66869 M25:GATE M25:DRN 2.943e-17
CC66855 M25:GATE M24:GATE 9.75e-18
R29 CP M11:GATE 125.306 
CC66851 CP N_42:1 2.397e-17
CC66817 CP N_42:1 8.584e-17
CC66882 CP M10:GATE 5.3e-18
CC66871 CP M25:DRN 4.53e-18
CC66894 CP M11:DRN 1.481e-17
CC66813 M11:GATE N_42:1 6.15e-18
CC66875 M11:GATE M10:GATE 9.95e-18
CC66872 M11:GATE M25:DRN 1e-18
CC66893 M11:GATE M11:DRN 2.325e-17
C30 M25:GATE 0 4.189e-17
C31 CP 0 1.926e-17
C32 M11:GATE 0 3.928e-17
R33 M1:GATE M22:SRC 240.775 
R34 M3:DRN M22:SRC 76.4371 
R35 M22:SRC M28:GATE 432.97 
CC66806 M22:SRC N_42:1 3.14e-17
CC67061 M22:SRC N_8:1 6.676e-17
CC66862 M22:SRC M22:GATE 1.468e-17
CC66843 M22:SRC N_42:1 1.74e-18
CC66821 M22:SRC N_42:2 2.702e-17
CC66737 M22:SRC M30:GATE 2.79e-17
CC66764 M22:SRC N_40:1 9.455e-17
CC66740 M22:SRC D 4.08e-18
CC66742 M22:SRC M3:GATE 1.94e-18
R36 M1:GATE M28:GATE 319.562 
R37 M28:GATE M3:DRN 417.899 
CC67063 M28:GATE N_8:1 7.93e-18
CC66845 M28:GATE N_42:1 4.38e-18
CC66911 M28:GATE M23:GATE 7.01e-18
CC66823 M28:GATE N_42:2 2.23e-18
CC67114 M28:GATE M28:SRC 2.105e-17
CC66765 M28:GATE N_40:1 4.061e-17
CC67103 M28:GATE M29:GATE 1.1e-18
R38 M3:DRN M1:GATE 232.391 
CC66798 M3:DRN M4:GATE 3.891e-17
CC66866 M3:DRN M22:GATE 7.26e-18
CC67134 M3:DRN M5:SRC 1e-18
CC66916 M3:DRN M8:GATE 1.733e-17
CC67076 M3:DRN N_8:1 2.64e-18
CC66800 M3:DRN M4:GATE 1.64e-18
CC66914 M3:DRN M23:GATE 5.73e-18
CC66830 M3:DRN N_42:2 1.55e-18
CC66771 M3:DRN N_40:1 8.43e-18
CC66735 M3:DRN M23:DRN 1.965e-17
CC66773 M3:DRN N_40:1 5.06e-18
CC66736 M3:DRN M22:DRN 1.912e-17
CC66741 M3:DRN D 9.495e-17
CC67126 M3:DRN M2:GATE 6.22e-18
CC67117 M3:DRN M28:SRC 1.404e-17
CC66739 M3:DRN M30:GATE 5.04e-18
CC66743 M3:DRN M3:GATE 4.46e-18
CC67078 M1:GATE N_8:1 6.126e-17
CC66910 M1:GATE CDN:2 1.07e-18
CC66774 M1:GATE N_40:1 1.85e-18
C39 M22:SRC 0 5.53e-18
C40 M28:GATE 0 4.054e-17
C41 M3:DRN 0 1.9e-17
C42 M1:GATE 0 2.3e-17
R43 M22:DRN M23:DRN 60.6736 
CC66822 M22:DRN N_42:2 2.48e-18
CC67123 M22:DRN M2:GATE 4.51e-18
CC66812 M22:DRN N_42:1 6.104e-17
CC67107 M22:DRN M29:GATE 2.305e-17
CC66913 M22:DRN M23:GATE 3.56e-18
CC67068 M22:DRN N_8:1 1.32e-18
CC66828 M22:DRN N_42:2 2.43e-18
CC66848 M22:DRN N_42:1 3.43e-18
CC66865 M22:DRN M22:GATE 3.415e-17
CC66912 M23:DRN M23:GATE 3.179e-17
CC67105 M23:DRN M29:GATE 3.421e-17
CC66811 M23:DRN N_42:1 1.21e-18
CC67067 M23:DRN N_8:1 5.751e-17
CC66827 M23:DRN N_42:2 4.45e-18
CC66915 M23:DRN M8:GATE 1.37e-18
C44 M22:DRN 0 1.542e-17
C45 M23:DRN 0 1.19e-17
R46 M3:GATE M30:GATE 531.699 
R47 M30:GATE D 142.349 
CC66783 M30:GATE M32:GATE 2.115e-17
CC66842 M30:GATE N_42:1 3.08e-18
CC66861 M30:GATE M22:GATE 3.79e-18
CC66820 M30:GATE N_42:2 3.24e-18
CC66805 M30:GATE N_42:1 2.01e-18
R48 D M3:GATE 124.105 
CC66776 D N_40:1 6.319e-17
CC66890 D M6:GATE 1.261e-17
CC66785 D M32:GATE 8.25e-18
CC66802 D M4:GATE 3.32e-18
CC66816 D N_42:1 1.848e-17
CC66880 M3:GATE M10:GATE 4.26e-18
CC66799 M3:GATE M4:GATE 2.12e-18
CC66772 M3:GATE N_40:1 2.383e-17
C49 M30:GATE 0 4.265e-17
C50 D 0 1.228e-17
C51 M3:GATE 0 2.643e-17
R52 M7:GATE M4:GATE 4532.81 
R53 M4:GATE N_40:1 87.6242 
CC67125 M4:GATE M2:GATE 1.571e-17
R54 M10:DRN N_40:1 30.2136 
R55 M32:GATE N_40:1 178.025 
R56 M24:DRN N_40:1 30.6279 
R57 M26:GATE N_40:1 262.306 
R58 N_40:1 M7:GATE 77.9282 
CC66818 N_40:1 N_42:1 1.123e-16
CC67127 N_40:1 M2:GATE 5.17e-18
CC67136 N_40:1 M5:SRC 1.034e-17
CC66895 N_40:1 M11:DRN 7.78e-18
CC66852 N_40:1 N_42:1 2.28e-18
CC66859 N_40:1 M24:GATE 9.38e-18
CC66883 N_40:1 M10:GATE 1.668e-17
CC66892 N_40:1 M6:GATE 5.45e-18
CC66970 N_40:1 M7:SRC 1.24e-18
CC66946 N_40:1 N_44:2 2.373e-17
CC67081 N_40:1 N_8:1 3.616e-17
CC66840 N_40:1 M9:GATE 5.89e-18
R59 M7:GATE M26:GATE 3764.08 
CC66833 M7:GATE M27:GATE 2.53e-18
CC67132 M7:GATE M5:SRC 2.076e-17
CC66969 M7:GATE M7:SRC 3.553e-17
CC66944 M7:GATE N_44:2 5.18e-18
CC67089 M7:GATE M27:DRN 2.08e-18
CC67073 M7:GATE N_8:1 5.83e-18
CC66838 M7:GATE M9:GATE 3.19e-18
CC66832 M26:GATE M27:GATE 2.01e-18
CC66937 M26:GATE N_44:2 8.5e-18
CC66951 M26:GATE M26:SRC 3.306e-17
CC66834 M26:GATE M9:GATE 5.96e-18
CC66810 M24:DRN N_42:1 1.445e-17
CC66856 M24:DRN M24:GATE 2.076e-17
CC66804 M32:GATE N_42:1 7.97e-18
CC66853 M32:GATE M24:GATE 1.01e-18
CC66873 M32:GATE M10:GATE 3.11e-18
CC66841 M32:GATE N_42:1 4.44e-18
CC66814 M10:DRN N_42:1 1.58e-18
CC66876 M10:DRN M10:GATE 3.66e-17
CC66887 M10:DRN M6:GATE 3.1e-18
C60 M4:GATE 0 2.454e-17
C61 N_40:1 0 3.8799e-16
C62 M7:GATE 0 1.03e-17
C63 M26:GATE 0 1.794e-17
C64 M24:DRN 0 1.816e-17
C65 M32:GATE 0 2.384e-17
C66 M10:DRN 0 1.664e-17
R67 M24:GATE N_42:1 165.97 
R68 N_42:2 N_42:1 1.31542 
R69 M11:DRN N_42:1 31.9685 
R70 M10:GATE N_42:1 131.252 
R71 N_42:1 M25:DRN 30.1961 
CC67110 N_42:1 M29:GATE 1.36e-18
CC67080 N_42:1 N_8:1 1.213e-17
CC67109 N_42:1 M29:GATE 5.5e-18
CC67118 N_42:1 M28:SRC 1.42e-18
R72 M6:GATE M10:GATE 248.041 
R73 M24:GATE M10:GATE 640.448 
R74 M10:GATE M11:DRN 5293.67 
R75 M22:GATE N_42:2 72.1458 
CC67106 M22:GATE M29:GATE 2.5e-18
R76 N_42:2 M27:GATE 81.0663 
CC67112 N_42:2 M29:GATE 5.51e-18
CC67121 N_42:2 M28:SRC 7.99e-18
CC67093 N_42:2 M27:DRN 2.913e-17
CC66947 N_42:2 N_44:2 2.704e-17
CC66955 N_42:2 M26:SRC 1.238e-17
CC67082 N_42:2 N_8:1 7.998e-17
R77 M27:GATE M9:GATE 134.941 
CC66950 M27:GATE M26:SRC 2.122e-17
CC66936 M27:GATE N_44:2 3.1e-18
CC66965 M27:GATE M7:SRC 1.097e-17
CC67086 M27:GATE M27:DRN 1.305e-17
CC67064 M27:GATE N_8:1 1.04e-18
CC66942 M9:GATE N_44:2 7.64e-18
CC66967 M9:GATE M7:SRC 2.352e-17
CC67070 M9:GATE N_8:1 1.3e-18
C78 N_42:1 0 2.7051e-16
C79 M25:DRN 0 1.465e-17
C80 M6:GATE 0 8.271e-17
C81 M10:GATE 0 7.986e-17
C82 M11:DRN 0 1.347e-17
C83 M22:GATE 0 1.414e-17
C84 N_42:2 0 1.2869e-16
C85 M27:GATE 0 2.8e-17
C86 M9:GATE 0 9.52e-18
C87 M24:GATE 0 1.339e-17
R88 M35:GATE CDN:1 154.043 
R89 M15:GATE CDN:1 119.715 
R90 CDN CDN:1 0.22 
R91 M18:GATE CDN:1 123.539 
R92 CDN:1 M38:GATE 149.235 
CC66993 CDN:1 N_15:1 7.568e-17
CC67005 CDN:1 M34:GATE 1.78e-18
CC66999 CDN:1 N_15:2 1.584e-17
CC66960 CDN:1 M16:GATE 1.024e-17
CC66935 CDN:1 M36:GATE 7.02e-18
CC66949 CDN:1 N_44:2 5.69e-17
CC66923 CDN:1 N_44:1 2.649e-17
CC66964 CDN:1 M17:GATE 3.72e-18
CC66929 CDN:1 M37:GATE 7.18e-18
CC67058 CDN:1 M16:SRC 1.127e-17
CC67043 CDN:1 M19:GATE 1.375e-17
CC67023 CDN:1 M35:SRC 1.33e-17
CC67016 CDN:1 M37:SRC 2.012e-17
CC67035 CDN:1 M21:GATE 1.002e-17
R93 M38:GATE M18:GATE 554.656 
CC66918 M38:GATE N_44:1 6.94e-18
CC66973 M38:GATE N_15:1 5.56e-18
CC67009 M38:GATE M37:SRC 9.73e-18
CC67025 M38:GATE M21:GATE 1.5e-18
R94 M18:GATE CDN:2 688.997 
CC66982 M18:GATE N_15:1 1.11e-18
CC66961 M18:GATE M17:GATE 3.52e-18
CC66940 M18:GATE N_44:2 4.61e-18
CC66920 M18:GATE N_44:1 9.41e-18
CC67037 M18:GATE M19:GATE 1.53e-18
R95 CDN:2 M8:GATE 109.975 
CC66972 CDN:2 M7:SRC 2.33e-18
CC66963 CDN:2 M17:GATE 5.45e-18
CC67138 CDN:2 M5:SRC 2.78e-18
CC67042 CDN:2 M19:GATE 3.17e-18
R96 M8:GATE M23:GATE 129.849 
CC67124 M8:GATE M2:GATE 5.59e-18
CC67072 M8:GATE N_8:1 7.84e-18
CC67104 M23:GATE M29:GATE 2.27e-18
CC67066 M23:GATE N_8:1 1.867e-17
CC66945 CDN N_44:2 4.102e-17
CC66922 CDN N_44:1 3.26e-18
CC66926 CDN M37:GATE 4.24e-18
CC67014 CDN M37:SRC 2.54e-18
R97 M15:GATE M35:GATE 522.444 
CC66985 M15:GATE N_15:1 2.97e-18
CC66996 M15:GATE N_15:2 2.283e-17
CC66957 M15:GATE M16:GATE 4.35e-18
CC67051 M15:GATE M14:GATE 3.38e-18
CC67002 M35:GATE M34:GATE 1.429e-17
CC66931 M35:GATE M36:GATE 6.46e-18
CC66976 M35:GATE N_15:1 2.589e-17
CC66919 M35:GATE N_44:1 2.7e-18
CC67020 M35:GATE M35:SRC 2.948e-17
C98 CDN:1 0 7.378e-17
C99 M38:GATE 0 3.468e-17
C100 M18:GATE 0 6.084e-17
C101 CDN:2 0 3.7279e-16
C102 M8:GATE 0 4.537e-17
C103 M23:GATE 0 2.596e-17
C104 CDN 0 1.1e-18
C105 M15:GATE 0 2.351e-17
C106 M35:GATE 0 2.969e-17
R107 M26:SRC N_44:2 29.9999 
R108 N_44:1 N_44:2 57.3028 
R109 M36:GATE N_44:2 278.83 
R110 M16:GATE N_44:2 235.934 
R111 N_44:2 M7:SRC 30.9024 
CC67095 N_44:2 M27:DRN 2.93e-18
CC67022 N_44:2 M35:SRC 2.04e-18
CC66992 N_44:2 N_15:1 1.4027e-16
CC67128 N_44:2 M2:GATE 4.75e-18
CC67015 N_44:2 M37:SRC 7.28e-18
CC67084 N_44:2 N_8:1 5.834e-17
CC67034 N_44:2 M21:GATE 5.27e-18
CC67057 N_44:2 M16:SRC 1.265e-17
CC67069 M7:SRC N_8:1 1.85e-18
CC67088 M7:SRC M27:DRN 1.19e-18
R112 N_44:1 M16:GATE 205.391 
R113 M16:GATE M36:GATE 999.41 
CC66984 M16:GATE N_15:1 5.47e-18
CC67055 M16:GATE M16:SRC 2.97e-18
R114 M36:GATE N_44:1 242.733 
CC67019 M36:GATE M35:SRC 2.944e-17
CC66975 M36:GATE N_15:1 6.71e-18
R115 M37:GATE N_44:1 104.675 
R116 N_44:1 M17:GATE 100.7 
CC67000 N_44:1 N_15:2 6.1e-18
CC67059 N_44:1 M16:SRC 4.492e-17
CC66983 M17:GATE N_15:1 3.12e-18
CC67054 M17:GATE M16:SRC 3.18e-18
CC67010 M37:GATE M37:SRC 2.918e-17
CC66974 M37:GATE N_15:1 6.99e-18
C117 M26:SRC 0 1.765e-17
C118 N_44:2 0 7.297e-17
C119 M7:SRC 0 5.38e-18
C120 M16:GATE 0 3.127e-17
C121 M36:GATE 0 3.527e-17
C122 N_44:1 0 2.096e-17
C123 M17:GATE 0 2.267e-17
C124 M37:GATE 0 2.436e-17
R125 M35:SRC M16:SRC 1784.09 
R126 N_15:1 M16:SRC 35.4755 
R127 M16:SRC N_15:2 498.612 
R128 M13:GATE N_15:2 144.124 
R129 M33:GATE N_15:2 170.513 
R130 M35:SRC N_15:2 1262.83 
R131 N_15:1 N_15:2 25.1107 
R132 M34:GATE N_15:2 111.3 
R133 N_15:2 M14:GATE 82.8124 
R134 M37:SRC N_15:1 29.9999 
R135 M35:SRC N_15:1 31.8903 
R136 N_15:1 M21:GATE 98.6578 
R137 M21:GATE M19:GATE 159 
R138 M33:GATE M13:GATE 591.409 
C139 M16:SRC 0 1.836e-17
C140 N_15:2 0 1.389e-17
C141 M14:GATE 0 1.832e-17
C142 M34:GATE 0 2.139e-17
C143 N_15:1 0 2.3373e-16
C144 M21:GATE 0 2.221e-17
C145 M19:GATE 0 3.551e-17
C146 M35:SRC 0 6.2e-18
C147 M33:GATE 0 3.064e-17
C148 M13:GATE 0 2.506e-17
C149 M37:SRC 0 6.02e-18
R150 M5:SRC N_8:1 30.4926 
R151 M28:SRC N_8:1 30.5038 
R152 M27:DRN N_8:1 30.3335 
R153 M29:GATE N_8:1 230.835 
R154 N_8:1 M2:GATE 86.6249 
R155 M2:GATE M29:GATE 528.598 
C156 M5:SRC 0 8.6e-19
C157 N_8:1 0 2.939e-17
C158 M2:GATE 0 6.74e-18
C159 M29:GATE 0 3.344e-17
C160 M27:DRN 0 1.166e-17
C161 M28:SRC 0 4.48e-18
.ENDS
*.SCALE METER 
.GLOBAL VSS VDD
