.SUBCKT BUFFD3 I Z
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.9e-07  AD=8e-14  AS=4.3e-14  PD=1.19e-06  PS=6.1e-07  SA=2.05e-07  SB=9.6e-07  NRD=0.648  NRS=1.112  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=9.95e-07  SB=1.6e-07  NRD=0.462  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.45e-07  SB=4.2e-07  NRD=4.183  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4.3e-14  PD=5.9e-07  PS=6.1e-07  SA=4.85e-07  SB=6.8e-07  NRD=4.141  NRS=1.112  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 M5:DRN M5:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=1.07e-13  AS=5.7e-14  PD=1.45e-06  PS=7.4e-07  SA=2.05e-07  SB=9.6e-07  NRD=0.569  NRS=0.293  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=9.95e-07  SB=1.6e-07  NRD=0.427  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vdd M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7.45e-07  SB=4.2e-07  NRD=2.057  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.7e-14  PD=7.2e-07  PS=7.4e-07  SA=4.85e-07  SB=6.8e-07  NRD=2.057  NRS=0.293  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M6:DRN Z 15.3824 
R1 M2:DRN Z 15.2993 
R2 M4:DRN Z 15.8699 
R3 Z M8:DRN 16.0118 
CC77823 Z M2:GATE 2.74e-18
CC77822 Z M6:GATE 1.127e-17
CC77801 Z N_6:1 3.387e-17
CC77810 Z M5:DRN 7.677e-17
CC77814 Z M8:GATE 5.52e-18
CC77807 Z N_6:2 3.47e-18
CC77819 Z M7:GATE 4.68e-18
CC77835 Z M1:DRN 1.97e-17
CC77826 Z M3:GATE 4.3e-18
CC77831 Z M4:GATE 2.71e-18
R4 M4:DRN M8:DRN 1025.82 
R5 M8:DRN M7:SRC 0.001 
CC77795 M8:DRN N_6:1 1.668e-17
CC77812 M8:DRN M8:GATE 4.577e-17
CC77816 M8:DRN M7:GATE 4.583e-17
CC77803 M8:DRN N_6:2 1.66e-18
R6 M4:DRN M3:SRC 0.001 
CC77798 M4:DRN N_6:1 5.506e-17
CC77805 M4:DRN N_6:2 4.14e-17
CC77833 M4:DRN M4:GATE 1.208e-17
CC77828 M4:DRN M3:GATE 8.68e-18
CC77825 M2:DRN M2:GATE 4.189e-17
CC77806 M2:DRN N_6:2 8.35e-18
CC77821 M6:DRN M6:GATE 4.589e-17
CC77804 M6:DRN N_6:2 1.66e-18
C7 Z 0 2.9132e-16
C8 M8:DRN 0 1.67e-17
C9 M4:DRN 0 8.57e-18
C10 M2:DRN 0 2.484e-17
C11 M6:DRN 0 2.588e-17
R12 M5:GATE M1:GATE 521.343 
R13 M1:GATE I 119.123 
CC77832 M1:GATE M4:GATE 1.59e-18
CC77800 M1:GATE N_6:1 1.56e-17
R14 I M5:GATE 145.077 
CC77830 I M4:GATE 2.68e-18
CC77836 I M1:DRN 3.69e-17
CC77815 I M8:GATE 1.74e-18
CC77802 I N_6:1 7.736e-17
CC77811 I M5:DRN 9.02e-18
CC77813 M5:GATE M8:GATE 5.94e-18
CC77834 M5:GATE M1:DRN 3.29e-18
CC77797 M5:GATE N_6:1 1.489e-17
CC77809 M5:GATE M5:DRN 2.783e-17
C15 M1:GATE 0 5.59e-17
C16 I 0 3.141e-17
C17 M5:GATE 0 7.858e-17
R18 M4:GATE N_6:1 81.2035 
R19 M8:GATE N_6:1 111.3 
R20 M5:DRN N_6:1 75.0338 
R21 M1:DRN N_6:1 74.8112 
R22 N_6:1 N_6:2 28.0588 
R23 M3:GATE N_6:2 94.0755 
R24 M7:GATE N_6:2 111.3 
R25 M6:GATE N_6:2 164.389 
R26 N_6:2 M2:GATE 138.947 
R27 M2:GATE M6:GATE 635.948 
R28 M1:DRN M5:DRN 105.307 
C29 N_6:1 0 8.362e-17
C30 N_6:2 0 4.592e-17
C31 M2:GATE 0 3.184e-17
C32 M6:GATE 0 1.007e-16
C33 M1:DRN 0 9.747e-17
C34 M5:DRN 0 4.524e-17
C35 M8:GATE 0 7.368e-17
C36 M7:GATE 0 9.363e-17
C37 M4:GATE 0 4.797e-17
C38 M3:GATE 0 5.052e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
