.SUBCKT INVD6 I ZN
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.9e-14  PD=7.2e-07  PS=7.1e-07  SA=6.7e-07  SB=9.3e-07  NRD=2.099  NRS=4.571  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.9e-14  AS=5.2e-14  PD=7.1e-07  PS=7.2e-07  SA=4.2e-07  SB=1.18e-06  NRD=4.571  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.567  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=1.44e-06  NRD=2.099  NRS=0.532  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.7e-14  PD=5.9e-07  PS=5.8e-07  SA=1.18e-06  SB=4.2e-07  NRD=4.141  NRS=6.091  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.7e-14  AS=3.9e-14  PD=5.8e-07  PS=5.9e-07  SA=9.3e-07  SB=6.7e-07  NRD=6.091  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.7e-14  PD=5.9e-07  PS=5.8e-07  SA=6.7e-07  SB=9.3e-07  NRD=4.141  NRS=6.091  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.7e-14  AS=3.9e-14  PD=5.8e-07  PS=5.9e-07  SA=4.2e-07  SB=1.18e-06  NRD=6.091  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.2e-14  PD=5.9e-07  PS=1.1e-06  SA=1.6e-07  SB=1.44e-06  NRD=4.141  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vdd M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.532  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.9e-14  PD=7.2e-07  PS=7.1e-07  SA=1.18e-06  SB=4.2e-07  NRD=2.099  NRS=4.571  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.9e-14  AS=5.2e-14  PD=7.1e-07  PS=7.2e-07  SA=9.3e-07  SB=6.7e-07  NRD=4.571  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M12:DRN M10:DRN 877.833 
R1 ZN M10:DRN 15.4615 
R2 M10:DRN M9:SRC 0.001 
CC38253 M10:DRN I:2 1.58e-18
CC38263 M10:DRN I:3 1.327e-17
CC38247 M10:DRN I:1 1.61e-18
CC38271 M10:DRN M9:GATE 4.576e-17
CC38269 M10:DRN M10:GATE 4.586e-17
R3 ZN M6:DRN 15.6009 
R4 M6:DRN M5:SRC 0.001 
CC38265 M6:DRN I:3 6.507e-17
CC38289 M6:DRN M5:GATE 8.24e-18
CC38286 M6:DRN M6:GATE 4.18e-17
CC38282 M6:DRN I 1.43e-18
R5 M2:DRN M4:DRN 1089.98 
R6 ZN M4:DRN 15.3877 
R7 M4:DRN M3:SRC 0.001 
CC38255 M4:DRN I:2 5.974e-17
CC38249 M4:DRN I:1 1.662e-17
CC38283 M4:DRN I 1.535e-17
CC38294 M4:DRN M3:GATE 1.406e-17
CC38293 M4:DRN M4:GATE 8.25e-18
R8 M2:DRN ZN 15.7222 
R9 M8:DRN ZN 15.7849 
R10 ZN M12:DRN 15.9342 
CC38256 ZN I:2 3.49e-18
CC38258 ZN M12:GATE 5.34e-18
CC38260 ZN M11:GATE 9.96e-18
CC38251 ZN I:1 5.77e-18
CC38291 ZN M4:GATE 8e-18
CC38288 ZN M5:GATE 4.5e-18
CC38287 ZN M6:GATE 1.601e-17
CC38285 ZN I 1.315e-16
CC38280 ZN M7:GATE 5.2e-18
CC38276 ZN M8:GATE 1.284e-17
CC38275 ZN M9:GATE 1.431e-17
CC38270 ZN M10:GATE 1.15e-17
CC38267 ZN I:3 4.31e-18
CC38300 ZN M1:GATE 3.8e-18
CC38297 ZN M2:GATE 8e-18
CC38296 ZN M3:GATE 6.71e-18
R11 M12:DRN M11:SRC 0.001 
CC38257 M12:DRN M12:GATE 4.605e-17
CC38259 M12:DRN M11:GATE 4.62e-17
CC38262 M12:DRN I:3 1.646e-17
CC38281 M12:DRN I 1.48e-18
R12 M8:DRN M7:SRC 0.001 
CC38264 M8:DRN I:3 1.331e-17
CC38248 M8:DRN I:1 3.33e-18
CC38279 M8:DRN M7:GATE 4.593e-17
CC38278 M8:DRN M8:GATE 4.582e-17
R13 M2:DRN M1:SRC 0.001 
CC38250 M2:DRN I:1 7.097e-17
CC38284 M2:DRN I 1.531e-17
CC38301 M2:DRN M1:GATE 2.024e-17
CC38299 M2:DRN M2:GATE 8.24e-18
C14 M10:DRN 0 6.58e-18
C15 M6:DRN 0 1.175e-17
C16 M4:DRN 0 7.26e-18
C17 ZN 0 3.4444e-16
C18 M12:DRN 0 1.051e-17
C19 M8:DRN 0 1.012e-17
C20 M2:DRN 0 1.116e-17
R21 I:2 I:3 22.9146 
R22 M11:GATE I:3 111.3 
R23 M5:GATE I:3 86.5669 
R24 M12:GATE I:3 269.655 
R25 M6:GATE I:3 200.636 
R26 I:3 I 16.0933 
R27 M12:GATE I 279.405 
R28 I M6:GATE 207.891 
R29 M6:GATE M12:GATE 1027.57 
R30 M10:GATE I:2 111.3 
R31 M4:GATE I:2 94.0755 
R32 M3:GATE I:2 236.785 
R33 M9:GATE I:2 280.141 
R34 I:2 I:1 58.8528 
R35 M8:GATE I:1 111.3 
R36 M2:GATE I:1 94.0755 
R37 M7:GATE I:1 164.389 
R38 M1:GATE I:1 138.947 
R39 M3:GATE I:1 227.678 
R40 I:1 M9:GATE 269.366 
R41 M9:GATE M3:GATE 1083.75 
R42 M1:GATE M7:GATE 635.948 
C43 I:3 0 4.859e-17
C44 I 0 1.0207e-16
C45 M6:GATE 0 2.721e-17
C46 M12:GATE 0 9.592e-17
C47 M5:GATE 0 4.171e-17
C48 M11:GATE 0 5.709e-17
C49 I:2 0 1.04e-18
C50 I:1 0 2.023e-17
C51 M9:GATE 0 4.825e-17
C52 M3:GATE 0 3.395e-17
C53 M4:GATE 0 3.468e-17
C54 M10:GATE 0 4.955e-17
C55 M1:GATE 0 6.16e-17
C56 M7:GATE 0 7.173e-17
C57 M2:GATE 0 4.167e-17
C58 M8:GATE 0 5.667e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
