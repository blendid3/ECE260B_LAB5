.SUBCKT INVD4 I ZN
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7e-14  AS=3.9e-14  PD=1.14e-06  PS=5.9e-07  SA=9.85e-07  SB=1.8e-07  NRD=0.508  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.25e-07  SB=4.4e-07  NRD=4.141  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.65e-07  SB=7e-07  NRD=4.183  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=8e-14  PD=5.9e-07  PS=1.19e-06  SA=2.05e-07  SB=9.6e-07  NRD=4.141  NRS=0.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=5.2e-07  AD=9.4e-14  AS=5.2e-14  PD=1.4e-06  PS=7.2e-07  SA=9.85e-07  SB=1.8e-07  NRD=0.453  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7.25e-07  SB=4.4e-07  NRD=2.057  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vdd M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.65e-07  SB=7e-07  NRD=2.099  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=1.07e-13  PD=7.2e-07  PS=1.45e-06  SA=2.05e-07  SB=9.6e-07  NRD=2.057  NRS=0.569  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M6:DRN ZN 15.614 
R1 M2:DRN ZN 15.5484 
R2 M4:DRN ZN 15.2802 
R3 ZN M8:DRN 15.338 
CC38222 ZN I:2 8.87e-18
CC38224 ZN M8:GATE 5.3e-18
CC38242 ZN M3:GATE 6.37e-18
CC38227 ZN M7:GATE 1.459e-17
CC38243 ZN M2:GATE 1.78e-18
CC38217 ZN I:1 2.101e-17
CC38238 ZN M4:GATE 2.82e-18
CC38237 ZN I 4.079e-17
CC38232 ZN M5:GATE 6.3e-18
CC38230 ZN M6:GATE 8.88e-18
CC38246 ZN M1:GATE 3.62e-18
R4 M6:DRN M8:DRN 1696.13 
R5 M8:DRN M7:SRC 0.001 
CC38223 M8:DRN M8:GATE 4.61e-17
CC38225 M8:DRN M7:GATE 4.755e-17
CC38233 M8:DRN I 6.02e-18
CC38213 M8:DRN I:1 9.33e-18
R6 M3:SRC M4:DRN 0.001 
CC38220 M4:DRN I:2 2.429e-17
CC38235 M4:DRN I 4.75e-18
CC38239 M4:DRN M4:GATE 4.208e-17
CC38240 M4:DRN M3:GATE 8.65e-18
CC38215 M4:DRN I:1 3.678e-17
R7 M2:DRN M1:SRC 0.001 
CC38221 M2:DRN I:2 3.734e-17
CC38216 M2:DRN I:1 1.075e-17
CC38236 M2:DRN I 4.52e-18
CC38245 M2:DRN M1:GATE 2.064e-17
CC38244 M2:DRN M2:GATE 4.173e-17
R8 M5:SRC M6:DRN 0.001 
CC38219 M6:DRN I:2 1.72e-18
CC38234 M6:DRN I 1.317e-17
CC38231 M6:DRN M5:GATE 4.591e-17
CC38229 M6:DRN M6:GATE 4.745e-17
C9 ZN 0 3.4299e-16
C10 M8:DRN 0 9.66e-18
C11 M4:DRN 0 1.114e-17
C12 M2:DRN 0 1.194e-17
C13 M6:DRN 0 1.083e-17
R14 M4:GATE I:1 94.0755 
R15 M3:GATE I:1 233.022 
R16 M7:GATE I:1 275.689 
R17 M8:GATE I:1 111.3 
R18 I I:1 41.1734 
R19 I:1 I:2 60.2341 
R20 M2:GATE I:2 94.0755 
R21 M6:GATE I:2 111.3 
R22 M3:GATE I:2 233.022 
R23 M7:GATE I:2 275.689 
R24 M5:GATE I:2 164.389 
R25 I:2 M1:GATE 138.947 
R26 M1:GATE M5:GATE 635.948 
R27 M7:GATE M3:GATE 1066.52 
C28 I:1 0 8.862e-17
C29 I:2 0 6.007e-17
C30 M1:GATE 0 6.135e-17
C31 M5:GATE 0 1.055e-16
C32 I 0 8.673e-17
C33 M8:GATE 0 7.213e-17
C34 M7:GATE 0 8.008e-17
C35 M3:GATE 0 6.502e-17
C36 M6:GATE 0 7.501e-17
C37 M2:GATE 0 2.542e-17
C38 M4:GATE 0 2.166e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
