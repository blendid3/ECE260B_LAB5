.SUBCKT XOR2D0 A1 A2 Z
MMM10 M9:DRN M10:GATE vdd vdd pch L=6e-08 W=2.15e-07  AD=2.2e-14  AS=3.7e-14  PD=4.11e-07  PS=7.06e-07  SA=1.5e-07  SB=4.35e-07  NRD=0.513  NRS=0.972  SCA=17.254  SCB=0.019  SCC=0.002 
MMM11 M11:DRN M11:GATE vdd vdd pch L=6e-08 W=2.67e-07  AD=4.3e-14  AS=4.6e-14  PD=8.5e-07  PS=8.74e-07  SA=1.65e-07  SB=1.72e-07  NRD=0.72  NRS=0.869  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=2.04e-07  AD=3.6e-14  AS=2.4e-14  PD=7.6e-07  PS=4.45e-07  SA=1.047e-06  SB=1.85e-07  NRD=0.996  NRS=0.844  SCA=15.333  SCB=0.018  SCC=0.002 
MMM12 M8:SRC M12:GATE M9:SRC vdd pch L=6e-08 W=2.68e-07  AD=5.7e-14  AS=4.2e-14  PD=8.1e-07  PS=7.45e-07  SA=1.45e-07  SB=2.2e-07  NRD=0.853  NRS=0.638  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=2.04e-07  AD=2.4e-14  AS=2e-14  PD=4.45e-07  PS=3.95e-07  SA=6.86e-07  SB=4.95e-07  NRD=0.844  NRS=8.262  SCA=15.333  SCB=0.018  SCC=0.002 
MMM3 M2:SRC M3:GATE M3:SRC vss nch L=6e-08 W=2e-07  AD=2e-14  AS=2.9e-14  PD=3.95e-07  PS=5.2e-07  SA=3.41e-07  SB=7.55e-07  NRD=8.262  NRS=0.774  SCA=15.333  SCB=0.018  SCC=0.002 
MMM4 M3:SRC M4:GATE M4:SRC vss nch L=6e-08 W=2.04e-07  AD=2.9e-14  AS=3e-14  PD=5.2e-07  PS=5.72e-07  SA=2.24e-07  SB=3.93e-07  NRD=0.774  NRS=0.813  SCA=9.037  SCB=0.011  SCC=0.000424 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=1.99e-07  AD=3.5e-14  AS=2.1e-14  PD=7.5e-07  PS=4.25e-07  SA=1.8e-07  SB=4.72e-07  NRD=0.972  NRS=5.674  SCA=14.747  SCB=0.017  SCC=0.001 
MMM6 M4:SRC M6:GATE vss vss nch L=6.2e-08 W=1.93e-07  AD=3e-14  AS=2e-14  PD=5.58e-07  PS=4.15e-07  SA=3.58e-07  SB=3.8e-07  NRD=0.833  NRS=4.081  SCA=18.359  SCB=0.02  SCC=0.002 
MMM7 M7:DRN M7:GATE vdd vdd pch L=6e-08 W=2.66e-07  AD=4.4e-14  AS=3.9e-14  PD=8.6e-07  PS=6.35e-07  SA=3e-07  SB=1.7e-07  NRD=0.737  NRS=0.78  SCA=6.877  SCB=0.008  SCC=0.0002134 
MMM8 vdd M8:GATE M8:SRC vdd pch L=6e-08 W=2.69e-07  AD=3.9e-14  AS=5.7e-14  PD=6.35e-07  PS=8.1e-07  SA=2.15e-07  SB=2.41e-07  NRD=0.78  NRS=0.853  SCA=15.255  SCB=0.017  SCC=0.002 
MMM9 M9:DRN M9:GATE M9:SRC vdd pch L=6e-08 W=2.63e-07  AD=2.7e-14  AS=4.2e-14  PD=5.09e-07  PS=7.45e-07  SA=2.99e-07  SB=1.75e-07  NRD=9.503  NRS=0.638  SCA=15.255  SCB=0.017  SCC=0.002 
R0 M1:DRN Z 30.2705 
CC79654 M1:DRN M1:GATE 3.198e-17
R1 Z M7:DRN 30.5658 
CC79569 Z A2 1.053e-17
CC79635 Z M7:GATE 1.164e-17
CC79655 Z M1:GATE 4.01e-18
CC79666 Z M3:SRC 6.625e-17
CC79632 M7:DRN M7:GATE 2.978e-17
CC79645 M7:DRN M9:SRC 1.47e-18
C2 M1:DRN 0 1.577e-17
C3 Z 0 8.746e-17
C4 M7:DRN 0 2.51e-17
R5 M8:GATE A2 114.653 
R6 A2 M2:GATE 99.7709 
CC79576 A2 M8:SRC 8.78e-18
CC79580 A2 M2:SRC 7.026e-17
CC79593 A2 M3:GATE 7.18e-18
CC79636 A2 M7:GATE 4.53e-18
CC79656 A2 M1:GATE 4.297e-17
R7 M2:GATE M8:GATE 305.528 
CC79579 M2:GATE M2:SRC 2.014e-17
CC79592 M2:GATE M3:GATE 3.52e-18
CC79653 M2:GATE M1:GATE 4.38e-18
CC79578 M8:GATE M2:SRC 4.69e-18
CC79574 M8:GATE M8:SRC 1.59e-17
CC79572 M8:GATE M8:SRC 2.24e-18
CC79631 M8:GATE M7:GATE 4.02e-18
CC79644 M8:GATE M9:SRC 2.102e-17
C8 A2 0 3.053e-17
C9 M2:GATE 0 2.962e-17
C10 M8:GATE 0 3.755e-17
R11 M3:GATE M9:GATE 249.631 
R12 M5:DRN M9:GATE 219.641 
R13 M9:GATE M11:DRN 212.288 
CC79687 M9:GATE M4:SRC 5.65e-18
CC79677 M9:GATE M9:DRN 3.107e-17
CC79658 M9:GATE M3:SRC 5.06e-18
CC79642 M9:GATE M9:SRC 5.278e-17
CC79602 M9:GATE M12:GATE 4.24e-18
CC79627 M9:GATE M9:SRC 1.047e-17
CC79619 M9:GATE M4:GATE 3.23e-18
CC79584 M9:GATE M10:GATE 3.04e-18
R14 M11:DRN M5:DRN 71.0844 
CC79684 M11:DRN M4:SRC 2.749e-17
CC79674 M11:DRN M9:DRN 7.31e-18
CC79640 M11:DRN M9:SRC 2.43e-18
CC79612 M11:DRN M5:GATE 1.407e-17
CC79596 M11:DRN M11:GATE 3.654e-17
CC79606 M11:DRN A1 7.55e-18
CC79600 M11:DRN M12:GATE 2.1e-18
CC79629 M11:DRN M7:GATE 3.099e-17
CC79625 M11:DRN M9:SRC 2.5e-18
CC79581 M11:DRN M10:GATE 7.11e-18
CC79583 M11:DRN M2:SRC 1.04e-18
CC79609 M5:DRN A1 6.978e-17
CC79616 M5:DRN M5:GATE 2.911e-17
CC79663 M3:GATE M3:SRC 3.454e-17
CC79589 M3:GATE M8:SRC 8.19e-18
CC79591 M3:GATE M2:SRC 4.434e-17
CC79604 M3:GATE M12:GATE 1.79e-18
CC79621 M3:GATE M4:GATE 2.8e-18
C15 M9:GATE 0 6.816e-17
C16 M11:DRN 0 6.15e-17
C17 M5:DRN 0 9.721e-17
C18 M3:GATE 0 7.57e-18
R19 M12:GATE M11:GATE 343.175 
CC79599 M12:GATE M8:SRC 2.34e-18
CC79623 M12:GATE M9:SRC 2.01e-18
CC79637 M12:GATE M9:SRC 1.94e-17
CC79603 M12:GATE M8:SRC 9.38e-18
R20 A1 M11:GATE 193.98 
R21 M11:GATE M5:GATE 580.47 
CC79597 M11:GATE M10:GATE 1.42e-18
CC79673 M11:GATE M9:DRN 1.42e-18
CC79624 M11:GATE M9:SRC 4.34e-18
CC79639 M11:GATE M9:SRC 7e-18
R22 M4:GATE M5:GATE 339.465 
R23 M5:GATE A1 99.069 
CC79617 M5:GATE M2:SRC 1.303e-17
CC79689 M5:GATE M4:SRC 3.3e-18
CC79613 M5:GATE M10:GATE 5.36e-18
CC79668 A1 M3:SRC 1.81e-18
CC79607 A1 M10:GATE 1.608e-17
CC79608 A1 M6:GATE 1.36e-18
CC79694 A1 M4:SRC 2.604e-17
CC79682 A1 M9:DRN 1.23e-18
CC79662 M4:GATE M3:SRC 2.549e-17
CC79622 M4:GATE M2:SRC 1.676e-17
CC79695 M4:GATE N_12:2 1.51e-18
CC79690 M4:GATE M4:SRC 1.938e-17
C24 M12:GATE 0 5.383e-17
C25 M11:GATE 0 1.4035e-16
C26 M5:GATE 0 1.1232e-16
C27 A1 0 7.347e-17
C28 M4:GATE 0 4.258e-17
R29 M10:GATE M6:GATE 137.8 
R30 M8:SRC M6:GATE 167.8 
R31 M6:GATE M2:SRC 164.303 
CC79688 M6:GATE M4:SRC 2.414e-17
CC79671 M6:GATE N_12:1 2.47e-18
CC79660 M6:GATE M3:SRC 5.767e-17
R32 M2:SRC M8:SRC 74.1832 
CC79681 M2:SRC M9:DRN 1.877e-17
CC79664 M2:SRC M3:SRC 2.768e-17
CC79648 M2:SRC M9:SRC 1.27e-18
CC79696 M2:SRC N_12:2 2.13e-18
CC79693 M2:SRC M4:SRC 6.13e-18
CC79643 M8:SRC M9:SRC 6.213e-17
CC79638 M8:SRC M9:SRC 2.58e-18
CC79685 M10:GATE M4:SRC 1.761e-17
CC79675 M10:GATE M9:DRN 3.084e-17
C33 M6:GATE 0 5.852e-17
C34 M2:SRC 0 6.31e-18
C35 M8:SRC 0 1.2569e-16
C36 M10:GATE 0 3.795e-17
R37 M9:SRC M3:SRC 75.585 
R38 M7:GATE M3:SRC 371.43 
R39 M1:GATE M3:SRC 276.478 
R40 N_13:2 M3:SRC 13.0339 
R41 M3:SRC N_13:1 14.1036 
R42 N_13:1 N_13:2 28.8227 
R43 M9:SRC M1:GATE 268.723 
R44 M1:GATE M7:GATE 317.149 
R45 M7:GATE M9:SRC 361.012 
CC79676 M9:SRC M9:DRN 6.398e-17
CC79686 M9:SRC M4:SRC 1.96e-18
C46 M3:SRC 0 4.708e-17
C47 N_13:1 0 1.39e-18
C48 M1:GATE 0 3.966e-17
C49 M7:GATE 0 5.376e-17
C50 M9:SRC 0 2.442e-17
R51 M9:DRN M4:SRC 60.4296 
R52 N_12:2 M4:SRC 15.2664 
R53 M4:SRC N_12:1 24.3625 
R54 N_12:1 N_12:2 13.4962 
C55 M4:SRC 0 2.362e-17
C56 N_12:1 0 1.4e-19
C57 M9:DRN 0 5.37e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
