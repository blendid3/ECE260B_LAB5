.SUBCKT BUFFD12 I Z
MMM20 M19:SRC M20:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=4.04e-06  NRD=2.057  NRS=0.427  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 vdd M21:GATE M21:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=4.04e-06  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=3.78e-06  SB=4.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 vdd M23:GATE M23:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=3.54e-06  SB=6.6e-07  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 M24:DRN M24:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.28e-06  SB=9.2e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM25 vdd M25:GATE M25:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.02e-06  SB=1.18e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM26 M26:DRN M26:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.76e-06  SB=1.44e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM27 vdd M27:GATE M27:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.5e-06  SB=1.7e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM28 M28:DRN M28:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.24e-06  SB=1.96e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM29 vdd M29:GATE M29:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.98e-06  SB=2.22e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.76e-06  SB=1.44e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.5e-06  SB=1.7e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.4e-07  SB=3.26e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.24e-06  SB=1.96e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M1:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=3.52e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.98e-06  SB=2.22e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=3.78e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.72e-06  SB=2.48e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M3:SRC M4:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.2e-14  PD=5.9e-07  PS=1.1e-06  SA=1.6e-07  SB=4.04e-06  NRD=4.141  NRS=0.462  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vss M15:GATE M15:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.46e-06  SB=2.74e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=4.04e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.2e-06  SB=3e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=3.78e-06  SB=4.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 M17:DRN M17:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.4e-07  SB=3.26e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=3.54e-06  SB=6.6e-07  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M17:DRN M18:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=3.52e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.28e-06  SB=9.2e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vdd M19:GATE M19:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=3.78e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.02e-06  SB=1.18e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM30 M30:DRN M30:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.72e-06  SB=2.48e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM31 vdd M31:GATE M31:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.46e-06  SB=2.74e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM32 M32:DRN M32:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.2e-06  SB=3e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M1:GATE M17:GATE 576.069 
R1 M17:GATE I:2 172.964 
CC29408 M17:GATE M1:DRN 3e-18
CC29355 M17:GATE M32:GATE 1.335e-17
CC29238 M17:GATE N_15:3 4.2e-18
CC29225 M17:GATE N_15:2 1.036e-17
CC29391 M17:GATE M17:DRN 4.874e-17
R2 M1:GATE I:2 146.196 
R3 M18:GATE I:2 111.3 
R4 M2:GATE I:2 80.8704 
R5 I:1 I:2 23.85 
R6 I:2 I 22.2149 
CC29394 I:2 M17:DRN 3.41e-18
CC29414 I:2 M1:DRN 6.298e-17
CC29235 I:2 N_15:2 1.62e-18
R7 I I:1 22 
CC29405 I M3:SRC 2.15e-18
CC29412 I M1:DRN 1.24e-18
CC29233 I N_15:2 1.0925e-16
R8 M19:GATE I:1 111.3 
R9 M4:GATE I:1 132.389 
R10 M20:GATE I:1 156.63 
R11 I:1 M3:GATE 81.5607 
CC29406 I:1 M3:SRC 5.69e-17
CC29393 I:1 M17:DRN 1.33e-17
CC29413 I:1 M1:DRN 1.431e-17
CC29234 I:1 N_15:2 2.89e-18
CC29385 I:1 M19:SRC 1.475e-17
CC29403 M3:GATE M3:SRC 1.04e-17
CC29230 M3:GATE N_15:2 5.67e-18
R12 M20:GATE M4:GATE 709.654 
CC29222 M20:GATE N_15:2 2.568e-17
CC29381 M20:GATE M19:SRC 5.071e-17
CC29402 M4:GATE M3:SRC 4.271e-17
CC29302 M4:GATE N_15:10 5.45e-18
CC29229 M4:GATE N_15:2 1.63e-18
CC29410 M2:GATE M1:DRN 1.127e-17
CC29231 M2:GATE N_15:2 6.32e-18
CC29224 M18:GATE N_15:2 1.216e-17
CC29390 M18:GATE M17:DRN 4.938e-17
CC29223 M19:GATE N_15:2 1.019e-17
CC29382 M19:GATE M19:SRC 4.912e-17
CC29411 M1:GATE M1:DRN 1.925e-17
CC29241 M1:GATE N_15:3 7.67e-18
CC29232 M1:GATE N_15:2 7.06e-18
CC29340 M1:GATE M16:GATE 3.67e-18
C13 M17:GATE 0 3.376e-17
C14 I:2 0 3.29e-18
C15 I 0 1.786e-17
C16 I:1 0 5.956e-17
C17 M3:GATE 0 3.308e-17
C18 M20:GATE 0 8.109e-17
C19 M4:GATE 0 4.369e-17
C20 M2:GATE 0 2.843e-17
C21 M18:GATE 0 2.776e-17
C22 M19:GATE 0 4.031e-17
C23 M1:GATE 0 2.524e-17
R24 M11:SRC M12:DRN 0.001 
R25 M12:DRN Z:1 14.9999 
CC29274 M12:DRN N_15:6 1.883e-17
CC29397 M12:DRN M12:GATE 1.005e-17
CC29373 M12:DRN M28:GATE 4.66e-18
CC29401 M12:DRN M11:GATE 1.22e-17
CC29298 M12:DRN N_15:10 6.384e-17
R26 M6:DRN Z:1 15.6563 
R27 M16:DRN Z:1 15.4749 
R28 M10:DRN Z:1 15.0394 
R29 M14:DRN Z:1 15.2851 
R30 M8:DRN Z:1 15.4714 
R31 Z:1 Z 0.10123 
CC29272 Z:1 N_15:5 3.06e-18
CC29249 Z:1 M26:GATE 5.69e-18
CC29375 Z:1 M28:GATE 1.59e-18
CC29338 Z:1 M16:GATE 4.6e-18
CC29337 Z:1 M5:GATE 3.78e-18
CC29380 Z:1 M27:GATE 6.27e-18
CC29331 Z:1 M6:GATE 1.347e-17
CC29328 Z:1 M7:GATE 1.439e-17
CC29325 Z:1 M8:GATE 1.546e-17
CC29322 Z:1 M9:GATE 1.414e-17
CC29321 Z:1 M10:GATE 1.442e-17
CC29351 Z:1 M15:GATE 1.414e-17
CC29345 Z:1 M14:GATE 1.543e-17
CC29369 Z:1 M29:GATE 1.79e-18
CC29342 Z:1 M13:GATE 1.109e-17
CC29288 Z:1 N_15:9 5.29e-18
CC29284 Z:1 N_15:8 4.71e-18
CC29280 Z:1 N_15:7 4.04e-18
CC29276 Z:1 N_15:6 5.21e-18
CC29398 Z:1 M12:GATE 1.461e-17
CC29317 Z:1 N_15:12 1.51e-18
CC29399 Z:1 M11:GATE 6.88e-18
CC29308 Z:1 N_15:11 2.25e-18
CC29307 Z:1 N_15:10 7.548e-17
CC29415 Z:1 M1:DRN 4.67e-18
CC29237 Z:1 N_15:2 1.1747e-16
CC29219 Z:1 N_15:1 1.0912e-16
R32 Z Z:2 0.104 
CC29303 Z N_15:10 2.33e-18
R33 M26:DRN Z:2 15.3984 
R34 M24:DRN Z:2 15.767 
R35 M30:DRN Z:2 15.4487 
R36 M32:DRN Z:2 15.6346 
R37 M22:DRN Z:2 15.9495 
R38 Z:2 M28:DRN 14.9999 
CC29267 Z:2 M21:GATE 4.42e-18
CC29252 Z:2 M25:GATE 1.763e-17
CC29248 Z:2 M26:GATE 1.645e-17
CC29264 Z:2 M22:GATE 1.681e-17
CC29260 Z:2 M23:GATE 1.836e-17
CC29256 Z:2 M24:GATE 1.772e-17
CC29379 Z:2 M27:GATE 1.474e-17
CC29395 Z:2 M17:DRN 7.77e-18
CC29356 Z:2 M32:GATE 4.92e-18
CC29360 Z:2 M31:GATE 1.667e-17
CC29364 Z:2 M30:GATE 1.859e-17
CC29368 Z:2 M29:GATE 1.477e-17
CC29374 Z:2 M28:GATE 1.45e-17
CC29306 Z:2 N_15:10 3.251e-17
CC29236 Z:2 N_15:2 7.892e-17
CC29218 Z:2 N_15:1 7.22e-17
R39 M28:DRN M27:SRC 0.001 
CC29376 M28:DRN M27:GATE 4.495e-17
CC29372 M28:DRN M28:GATE 4.52e-17
CC29291 M28:DRN N_15:10 1.146e-17
R40 M24:DRN M22:DRN 753.317 
R41 M22:DRN M21:SRC 0.001 
CC29266 M22:DRN M21:GATE 4.626e-17
CC29263 M22:DRN M22:GATE 4.481e-17
CC29294 M22:DRN N_15:10 1.149e-17
CC29214 M22:DRN N_15:1 1.26e-18
R42 M6:DRN M8:DRN 990.169 
R43 M8:DRN M7:SRC 0.001 
CC29329 M8:DRN M7:GATE 5.07e-18
CC29326 M8:DRN M8:GATE 4.89e-18
CC29281 M8:DRN N_15:8 4.178e-17
CC29279 M8:DRN N_15:7 4.176e-17
CC29300 M8:DRN N_15:10 1.457e-17
CC29216 M8:DRN N_15:1 1.17e-18
R44 M31:SRC M32:DRN 0.001 
R45 M32:DRN M30:DRN 1039.16 
CC29357 M32:DRN M31:GATE 4.529e-17
CC29352 M32:DRN M32:GATE 4.646e-17
CC29289 M32:DRN N_15:10 1.154e-17
CC29220 M32:DRN N_15:2 1.44e-18
R46 M30:DRN M29:SRC 0.001 
CC29363 M30:DRN M30:GATE 4.597e-17
CC29366 M30:DRN M29:GATE 4.587e-17
CC29290 M30:DRN N_15:10 1.164e-17
CC29221 M30:DRN N_15:2 1.31e-18
R47 M16:DRN M14:DRN 1619.1 
R48 M14:DRN M13:SRC 0.001 
CC29273 M14:DRN N_15:6 4.259e-17
CC29347 M14:DRN M14:GATE 5.07e-18
CC29344 M14:DRN M13:GATE 5.07e-18
CC29311 M14:DRN N_15:11 4.22e-17
CC29297 M14:DRN N_15:10 1.457e-17
CC29227 M14:DRN N_15:2 1.5e-18
R49 M10:DRN M9:SRC 0.001 
CC29269 M10:DRN N_15:5 6.33e-17
CC29324 M10:DRN M9:GATE 6.39e-18
CC29320 M10:DRN M10:GATE 1.352e-17
CC29299 M10:DRN N_15:10 2.563e-17
R50 M26:DRN M24:DRN 878.324 
R51 M24:DRN M23:SRC 0.001 
CC29255 M24:DRN M24:GATE 4.51e-17
CC29258 M24:DRN M23:GATE 4.505e-17
CC29293 M24:DRN N_15:10 1.164e-17
CC29213 M24:DRN N_15:1 1.31e-18
R52 M26:DRN M25:SRC 0.001 
CC29250 M26:DRN M25:GATE 4.514e-17
CC29247 M26:DRN M26:GATE 4.495e-17
CC29292 M26:DRN N_15:10 1.16e-17
CC29212 M26:DRN N_15:1 1.03e-18
R53 M16:DRN M15:SRC 0.001 
CC29239 M16:DRN N_15:3 3.441e-17
CC29348 M16:DRN M15:GATE 6.39e-18
CC29341 M16:DRN M16:GATE 1.393e-17
CC29313 M16:DRN N_15:12 4.104e-17
CC29296 M16:DRN N_15:10 1.387e-17
CC29226 M16:DRN N_15:2 1.89e-18
R54 M6:DRN M5:SRC 0.001 
CC29335 M6:DRN M5:GATE 5.33e-18
CC29333 M6:DRN M6:GATE 5.1e-18
CC29286 M6:DRN N_15:9 5.865e-17
CC29301 M6:DRN N_15:10 1.378e-17
CC29217 M6:DRN N_15:1 2.712e-17
C55 M12:DRN 0 4.62e-18
C56 Z:1 0 2.7012e-16
C57 Z 0 5.9e-19
C58 Z:2 0 2.9503e-16
C59 M28:DRN 0 4.98e-18
C60 M22:DRN 0 1.882e-17
C61 M8:DRN 0 4e-18
C62 M32:DRN 0 8.05e-18
C63 M30:DRN 0 4.81e-18
C64 M14:DRN 0 4.62e-18
C65 M10:DRN 0 6.21e-18
C66 M24:DRN 0 1.584e-17
C67 M26:DRN 0 6.61e-18
C68 M16:DRN 0 4.85e-18
C69 M6:DRN 0 7.6e-18
R70 N_15:6 M12:GATE 259.951 
R71 N_15:10 M12:GATE 237.148 
R72 M12:GATE M28:GATE 1033.72 
R73 N_15:6 M28:GATE 277.281 
R74 M28:GATE N_15:10 252.958 
R75 M27:GATE N_15:10 83.475 
R76 N_15:6 N_15:10 63.6118 
R77 M11:GATE N_15:10 99.3746 
R78 N_15:5 N_15:10 59.4752 
R79 M26:GATE N_15:10 264.336 
R80 N_15:10 M10:GATE 247.815 
R81 N_15:5 M10:GATE 243.049 
R82 M10:GATE M26:GATE 1080.21 
R83 M26:GATE N_15:5 259.25 
R84 M25:GATE N_15:5 106 
R85 N_15:7 N_15:5 21.9882 
R86 M9:GATE N_15:5 91.8666 
R87 N_15:5 N_15:1 23.1924 
R88 N_15:7 N_15:1 23.1924 
R89 N_15:8 N_15:1 22.7027 
R90 M21:GATE N_15:1 322.403 
R91 M5:GATE N_15:1 302.252 
R92 N_15:1 N_15:9 15.0611 
R93 M22:GATE N_15:9 106 
R94 M6:GATE N_15:9 85.86 
R95 N_15:8 N_15:9 21.9794 
R96 M21:GATE N_15:9 271.188 
R97 N_15:9 M5:GATE 254.238 
R98 M5:GATE M21:GATE 732.576 
R99 M16:GATE N_15:3 87.2465 
R100 M32:GATE N_15:3 93.8715 
R101 N_15:12 N_15:3 22.8364 
R102 N_15:3 N_15:2 22.2205 
R103 N_15:6 N_15:2 22.2385 
R104 N_15:11 N_15:2 22 
R105 M19:SRC N_15:2 16.6394 
R106 M17:DRN N_15:2 16.0859 
R107 M1:DRN N_15:2 15.9398 
R108 M3:SRC N_15:2 16.4689 
R109 N_15:2 N_15:12 22.2294 
R110 M31:GATE N_15:12 96.9899 
R111 N_15:11 N_15:12 21.9794 
R112 N_15:12 M15:GATE 90.365 
R113 M3:SRC M1:DRN 546.12 
R114 M17:DRN M19:SRC 481.651 
R115 M7:GATE N_15:8 86.5037 
R116 M23:GATE N_15:8 106 
R117 N_15:8 N_15:7 22.6719 
R118 M24:GATE N_15:7 106 
R119 N_15:7 M8:GATE 89.1364 
R120 M14:GATE N_15:11 91.8666 
R121 N_15:6 N_15:11 22.4472 
R122 N_15:11 M30:GATE 98.4912 
R123 M29:GATE N_15:6 95.7611 
R124 N_15:6 M13:GATE 89.1364 
C125 M12:GATE 0 3.108e-17
C126 M28:GATE 0 4.743e-17
C127 N_15:10 0 1.0098e-16
C128 M10:GATE 0 2.179e-17
C129 M26:GATE 0 2.874e-17
C130 N_15:5 0 5.23e-18
C131 N_15:1 0 2.825e-17
C132 N_15:9 0 1.072e-17
C133 M5:GATE 0 6.566e-17
C134 M21:GATE 0 7.792e-17
C135 N_15:3 0 1.27e-18
C136 N_15:2 0 2.2679e-16
C137 N_15:12 0 2.29e-18
C138 M15:GATE 0 2.345e-17
C139 M11:GATE 0 3.553e-17
C140 M3:SRC 0 1.677e-17
C141 M1:DRN 0 7.55e-18
C142 M17:DRN 0 7.71e-18
C143 M19:SRC 0 2.35e-17
C144 M9:GATE 0 2.239e-17
C145 M7:GATE 0 2.408e-17
C146 N_15:8 0 4.61e-18
C147 N_15:7 0 7.89e-18
C148 M8:GATE 0 2.916e-17
C149 N_15:11 0 6.77e-18
C150 M30:GATE 0 5.078e-17
C151 N_15:6 0 1.97e-18
C152 M13:GATE 0 2.934e-17
C153 M6:GATE 0 3.231e-17
C154 M29:GATE 0 4.459e-17
C155 M27:GATE 0 4.862e-17
C156 M32:GATE 0 2.968e-17
C157 M31:GATE 0 3.447e-17
C158 M16:GATE 0 1.906e-17
C159 M14:GATE 0 3.323e-17
C160 M25:GATE 0 2.829e-17
C161 M24:GATE 0 2.165e-17
C162 M23:GATE 0 1.736e-17
C163 M22:GATE 0 2.403e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
