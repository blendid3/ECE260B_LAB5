.SUBCKT XOR2D1 A1 A2 Z
MMM10 vdd M10:GATE M10:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.4e-14  PD=7.2e-07  PS=1.004e-06  SA=3.55e-07  SB=4.35e-07  NRD=2.099  NRS=0.379  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 M7:SRC M11:GATE M10:SRC vdd pch L=6e-08 W=3.47e-07  AD=4.9e-14  AS=5.5e-14  PD=8e-07  PS=6.56e-07  SA=1.89e-07  SB=6.73e-07  NRD=0.459  NRS=0.503  SCA=4.486  SCB=0.003  SCC=4.492e-05 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.9e-07  AD=6.8e-14  AS=3.9e-14  PD=1.13e-06  PS=5.9e-07  SA=7.81e-07  SB=1.75e-07  NRD=0.496  NRS=4.183  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=2.67e-07  AD=4.3e-14  AS=4.6e-14  PD=8.5e-07  PS=8.74e-07  SA=1.65e-07  SB=1.72e-07  NRD=0.72  NRS=0.869  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4.1e-14  PD=5.9e-07  PS=6.48e-07  SA=4.25e-07  SB=4.35e-07  NRD=4.183  NRS=5.861  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM3 M2:SRC M3:GATE M3:SRC vss nch L=6e-08 W=3.28e-07  AD=3.3e-14  AS=4.3e-14  PD=5.32e-07  PS=6.45e-07  SA=3.73e-07  SB=6.95e-07  NRD=0.366  NRS=0.46  SCA=11.685  SCB=0.013  SCC=0.000978 
MMM4 M3:SRC M4:GATE M4:SRC vss nch L=6e-08 W=3.19e-07  AD=4.2e-14  AS=4.6e-14  PD=6.25e-07  PS=8.43e-07  SA=1.78e-07  SB=5.17e-07  NRD=0.471  NRS=0.521  SCA=7.393  SCB=0.008  SCC=0.0002747 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=1.99e-07  AD=3.5e-14  AS=2.1e-14  PD=7.5e-07  PS=4.25e-07  SA=1.8e-07  SB=4.72e-07  NRD=0.972  NRS=5.674  SCA=14.747  SCB=0.017  SCC=0.001 
MMM6 M4:SRC M6:GATE vss vss nch L=6.2e-08 W=1.93e-07  AD=2.8e-14  AS=2e-14  PD=5.17e-07  PS=4.15e-07  SA=3.58e-07  SB=3.78e-07  NRD=0.799  NRS=4.081  SCA=18.359  SCB=0.02  SCC=0.002 
MMM7 M7:DRN M7:GATE M7:SRC vdd pch L=6e-08 W=3.13e-07  AD=3.3e-14  AS=4.4e-14  PD=6.08e-07  PS=7.3e-07  SA=2.51e-07  SB=2.58e-07  NRD=11.086  NRS=0.493  SCA=13.685  SCB=0.015  SCC=0.001 
MMM8 M7:DRN M8:GATE vdd vdd pch L=6e-08 W=2.16e-07  AD=2.2e-14  AS=3.7e-14  PD=4.12e-07  PS=7.06e-07  SA=1.5e-07  SB=4.5e-07  NRD=0.523  NRS=0.972  SCA=17.254  SCB=0.019  SCC=0.002 
MMM9 M9:DRN M9:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=9.1e-14  AS=5.2e-14  PD=1.39e-06  PS=7.2e-07  SA=6.49e-07  SB=1.75e-07  NRD=0.541  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M9:DRN Z 30.6365 
CC80174 M9:DRN M9:GATE 2.902e-17
CC80187 M9:DRN M7:SRC 3.16e-18
R1 Z M1:DRN 15.2852 
CC80177 Z M9:GATE 1.309e-17
CC80222 Z M3:SRC 7.452e-17
CC80114 Z A2 1.218e-17
CC80206 Z M1:GATE 4.11e-18
CC80176 M1:DRN M9:GATE 7.27e-18
CC80221 M1:DRN M3:SRC 3.296e-17
CC80205 M1:DRN M1:GATE 1.353e-17
C2 M9:DRN 0 3.37e-17
C3 Z 0 1.1983e-16
C4 M1:DRN 0 2.448e-17
R5 M10:GATE M2:GATE 577.95 
R6 M2:GATE A2 124.874 
CC80196 M2:GATE M7:SRC 3.23e-18
CC80204 M2:GATE M1:GATE 3.66e-18
CC80115 M2:GATE M7:GATE 2.69e-18
CC80116 M2:GATE M3:GATE 2.86e-18
CC80117 M2:GATE M2:SRC 3.92e-18
R7 A2 M10:GATE 150.302 
CC80207 A2 M1:GATE 3.15e-18
CC80108 A2 M10:SRC 8.81e-18
CC80110 A2 M7:GATE 1.45e-18
CC80111 A2 M3:GATE 7.66e-18
CC80112 A2 M2:SRC 8.883e-17
CC80178 A2 M9:GATE 4.418e-17
CC80200 M10:GATE M1:GATE 6.72e-18
CC80103 M10:GATE M10:SRC 1.23e-17
CC80105 M10:GATE M2:SRC 5.06e-18
CC80186 M10:GATE M7:SRC 1.238e-17
CC80173 M10:GATE M9:GATE 7.1e-18
C8 M2:GATE 0 6.271e-17
C9 A2 0 4.101e-17
C10 M10:GATE 0 9.335e-17
R11 M11:GATE M12:GATE 348.476 
R12 M5:GATE M12:GATE 580.47 
R13 M12:GATE A1 193.98 
CC80128 M12:GATE M8:GATE 1.45e-18
CC80127 M12:GATE M12:DRN 3.662e-17
CC80182 M12:GATE M7:SRC 6.38e-18
CC80179 M12:GATE M7:SRC 3.71e-18
CC80149 M12:GATE M7:DRN 1.63e-18
R14 A1 M5:GATE 99.069 
CC80131 A1 M8:GATE 1.702e-17
CC80130 A1 M12:DRN 7.54e-18
CC80134 A1 M5:DRN 7.426e-17
CC80198 A1 M7:SRC 1.81e-18
CC80168 A1 M4:SRC 2.362e-17
CC80157 A1 M7:DRN 1.21e-18
R15 M5:GATE M4:GATE 332.045 
CC80165 M5:GATE M4:SRC 5.69e-18
CC80136 M5:GATE M12:DRN 1.406e-17
CC80137 M5:GATE M8:GATE 5e-18
CC80138 M5:GATE M6:GATE 1.237e-17
CC80139 M5:GATE M5:DRN 2.463e-17
CC80140 M5:GATE M2:SRC 2.02e-18
CC80218 M4:GATE M3:SRC 1.912e-17
CC80193 M4:GATE M7:SRC 6.84e-18
CC80166 M4:GATE M4:SRC 1.685e-17
CC80159 M4:GATE M4:SRC 4.54e-18
CC80142 M4:GATE M7:GATE 4.11e-18
CC80144 M4:GATE M3:GATE 3.75e-18
CC80145 M4:GATE M2:SRC 1.384e-17
CC80147 M4:GATE N_13:1 2.2e-18
CC80126 M11:GATE N_15:1 1.12e-18
CC80125 M11:GATE M2:SRC 1.25e-18
CC80124 M11:GATE M3:GATE 2.65e-18
CC80123 M11:GATE M7:GATE 4.29e-18
CC80121 M11:GATE M10:SRC 1.27e-17
CC80120 M11:GATE M12:DRN 2.2e-18
CC80185 M11:GATE M7:SRC 2.755e-17
C16 M12:GATE 0 1.4778e-16
C17 A1 0 7.098e-17
C18 M5:GATE 0 1.1522e-16
C19 M4:GATE 0 4.345e-17
C20 M11:GATE 0 4.328e-17
R21 M6:GATE M2:SRC 164.106 
R22 M2:SRC M10:SRC 74.2471 
CC80148 M2:SRC N_13:1 7.03e-18
CC80203 M2:SRC M1:GATE 1.207e-17
CC80210 M2:SRC M3:SRC 1.19e-18
CC80099 M2:SRC M3:GATE 3.611e-17
CC80175 M2:SRC M9:GATE 1.72e-18
CC80167 M2:SRC M4:SRC 1.692e-17
CC80195 M2:SRC M7:SRC 3.07e-18
CC80156 M2:SRC M7:DRN 1.879e-17
CC80220 M2:SRC M3:SRC 4.4e-18
CC80096 M2:SRC M7:GATE 1.246e-17
CC80092 M2:SRC M12:DRN 1.04e-18
R23 N_15:1 M10:SRC 10.7803 
R24 M10:SRC M6:GATE 167.794 
CC80184 M10:SRC M7:SRC 5.593e-17
CC80097 M10:SRC M3:GATE 8.19e-18
R25 M6:GATE M8:GATE 137.8 
CC80164 M6:GATE M4:SRC 1.764e-17
CC80216 M6:GATE M3:SRC 7.456e-17
CC80152 M8:GATE M7:DRN 3.259e-17
CC80162 M8:GATE M4:SRC 1.741e-17
CC80091 M8:GATE M12:DRN 6.7e-18
CC80094 M8:GATE M7:GATE 4.34e-18
C26 M2:SRC 0 5.16e-18
C27 M10:SRC 0 1.3545e-16
C28 M6:GATE 0 1.487e-17
C29 M8:GATE 0 3.634e-17
C30 N_15:1 0 1.01e-18
R31 M3:GATE M7:GATE 272.951 
CC80169 M3:GATE N_14:1 1.68e-18
CC80208 M3:GATE M3:SRC 1.2e-18
CC80194 M3:GATE M7:SRC 1.829e-17
CC80219 M3:GATE M3:SRC 2.39e-17
R32 M12:DRN M7:GATE 199.261 
R33 M7:GATE M5:DRN 206.16 
CC80181 M7:GATE M7:SRC 5.39e-18
CC80153 M7:GATE M7:DRN 3.195e-17
CC80163 M7:GATE M4:SRC 6.13e-18
CC80190 M7:GATE M7:SRC 3.959e-17
CC80215 M7:GATE M3:SRC 1.168e-17
R34 M5:DRN M12:DRN 71.8577 
CC80191 M5:DRN M7:SRC 2.99e-18
CC80150 M12:DRN M7:DRN 7.12e-18
CC80183 M12:DRN M7:SRC 2.93e-18
CC80161 M12:DRN M4:SRC 2.747e-17
CC80199 M12:DRN M1:GATE 3.079e-17
C35 M3:GATE 0 2.129e-17
C36 M7:GATE 0 6.812e-17
C37 M5:DRN 0 9.182e-17
C38 M12:DRN 0 6.154e-17
R39 M7:DRN M4:SRC 60.4296 
R40 M4:SRC N_13:1 10.6529 
CC80192 M4:SRC M7:SRC 2.07e-18
CC80189 M7:DRN M7:SRC 6.419e-17
C41 M4:SRC 0 2.147e-17
C42 N_13:1 0 1.1e-19
C43 M7:DRN 0 6.78e-18
R44 M3:SRC M9:GATE 345.821 
R45 M1:GATE M9:GATE 407.866 
R46 M9:GATE M7:SRC 336.121 
R47 M3:SRC M7:SRC 73.978 
R48 M7:SRC M1:GATE 340.935 
R49 M1:GATE M3:SRC 350.773 
R50 N_14:2 M3:SRC 30.0617 
R51 M3:SRC N_14:1 28.887 
R52 N_14:1 N_14:2 14.1489 
C53 M9:GATE 0 5.608e-17
C54 M7:SRC 0 4.12e-17
C55 M1:GATE 0 5.893e-17
C56 M3:SRC 0 4.696e-17
C57 N_14:1 0 2.3e-19
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
