.SUBCKT OR2D2 A1 A2 Z
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=2e-07  AD=3.7e-14  AS=2e-14  PD=7.7e-07  PS=4.05e-07  SA=1.9e-07  SB=1.015e-06  NRD=1.509  NRS=5.196  SCA=18.109  SCB=0.02  SCC=0.002 
MMM2 M1:SRC M2:GATE vss vss nch L=6e-08 W=2.04e-07  AD=2e-14  AS=2.9e-14  PD=4.05e-07  PS=4.27e-07  SA=4.6e-07  SB=7.45e-07  NRD=5.196  NRS=0.882  SCA=18.109  SCB=0.02  SCC=0.002 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=6.8e-14  AS=3.9e-14  PD=1.13e-06  PS=5.9e-07  SA=6.4e-07  SB=1.75e-07  NRD=0.592  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=5.8e-14  PD=5.9e-07  PS=8.53e-07  SA=3.27e-07  SB=4.35e-07  NRD=4.141  NRS=0.755  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 M5:DRN M5:GATE M5:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.6e-14  AS=5.5e-14  PD=1.37e-06  PS=7.3e-07  SA=1.65e-07  SB=1.035e-06  NRD=0.534  NRS=0.202  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M5:SRC M6:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.5e-14  AS=6.6e-14  PD=7.3e-07  PS=7.75e-07  SA=4.35e-07  SB=7.65e-07  NRD=0.202  NRS=0.657  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vdd M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=9.6e-14  AS=5.3e-14  PD=1.41e-06  PS=7.25e-07  SA=1.015e-06  SB=1.85e-07  NRD=0.549  NRS=1.051  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.3e-14  AS=6.6e-14  PD=7.25e-07  PS=7.75e-07  SA=7.5e-07  SB=4.5e-07  NRD=1.051  NRS=0.657  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 A1 M1:GATE 86.2084 
R1 M1:GATE M5:GATE 373.703 
CC11182 M1:GATE A2 4.03e-18
CC11181 M1:GATE M2:GATE 1.99e-18
CC11204 M1:GATE M5:DRN 1.52e-18
CC11213 M1:GATE M1:SRC 8.84e-18
CC11190 M1:GATE N_8:1 2.72e-18
R2 M5:GATE A1 157.582 
CC11177 M5:GATE A2 2.55e-18
CC11176 M5:GATE M6:GATE 1.259e-17
CC11203 M5:GATE M5:DRN 2.879e-17
CC11187 M5:GATE N_8:1 9.68e-18
CC11180 A1 A2 2.135e-17
CC11179 A1 M2:GATE 1.264e-17
CC11206 A1 M5:DRN 6.79e-18
CC11215 A1 M1:SRC 6.832e-17
C3 M1:GATE 0 4.584e-17
C4 M5:GATE 0 4.497e-17
C5 A1 0 4.18e-17
R6 A2 M2:GATE 88.872 
R7 M2:GATE M6:GATE 395.013 
CC11189 M2:GATE N_8:1 8.78e-18
CC11212 M2:GATE M1:SRC 8.79e-18
R8 M6:GATE A2 159.193 
CC11186 M6:GATE N_8:1 2.219e-17
CC11195 M6:GATE M8:GATE 4.66e-18
CC11214 A2 M1:SRC 2.749e-17
CC11201 A2 M7:GATE 1.64e-18
CC11207 A2 M4:GATE 2.32e-18
CC11198 A2 M8:GATE 1.54e-18
CC11205 A2 M5:DRN 8.685e-17
CC11192 A2 N_8:1 1.83e-18
C9 M2:GATE 0 3.187e-17
C10 M6:GATE 0 7.148e-17
C11 A2 0 1.416e-17
R12 M7:SRC M8:DRN 0.001 
R13 M8:DRN Z 15.5946 
CC11185 M8:DRN N_8:1 1.297e-17
CC11194 M8:DRN M8:GATE 4.249e-17
CC11199 M8:DRN M7:GATE 5.203e-17
R14 Z M4:DRN 15.2637 
CC11191 Z N_8:1 1.0508e-16
CC11197 Z M8:GATE 4.01e-18
CC11200 Z M7:GATE 1.58e-17
CC11208 Z M4:GATE 3.05e-18
CC11210 Z M3:GATE 1.26e-17
R15 M4:DRN M3:SRC 0.001 
CC11188 M4:DRN N_8:1 9.979e-17
CC11211 M4:DRN M3:GATE 7.49e-18
CC11209 M4:DRN M4:GATE 7.09e-18
C16 M8:DRN 0 1.074e-17
C17 Z 0 1.3698e-16
C18 M4:DRN 0 8.69e-18
R19 M8:GATE N_8:1 111.3 
R20 M1:SRC N_8:1 74.3102 
R21 M5:DRN N_8:1 76.0505 
R22 M4:GATE N_8:1 80.5597 
R23 M3:GATE N_8:1 139.81 
R24 N_8:1 M7:GATE 165.41 
R25 M7:GATE M3:GATE 627.823 
R26 M5:DRN M1:SRC 106.518 
C27 M8:GATE 0 6.71e-17
C28 N_8:1 0 5.537e-17
C29 M7:GATE 0 8.021e-17
C30 M3:GATE 0 7.072e-17
C31 M4:GATE 0 4.711e-17
C32 M5:DRN 0 6.43e-17
C33 M1:SRC 0 8.155e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
