.SUBCKT ND2D2 A1 A2 ZN
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=8e-14  AS=3.9e-14  PD=1.19e-06  PS=5.9e-07  SA=9.85e-07  SB=2.05e-07  NRD=0.566  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M1:SRC M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.25e-07  SB=4.65e-07  NRD=4.12  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.65e-07  SB=7.25e-07  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M3:SRC M4:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=8e-14  PD=5.9e-07  PS=1.19e-06  SA=2.05e-07  SB=9.85e-07  NRD=4.12  NRS=0.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=5.24e-07  AD=9.9e-14  AS=5.2e-14  PD=1.42e-06  PS=7.2e-07  SA=9.7e-07  SB=1.9e-07  NRD=1.471  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7.1e-07  SB=4.5e-07  NRD=2.099  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vdd M7:GATE M7:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.5e-07  SB=7.1e-07  NRD=2.534  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=9.9e-14  PD=7.2e-07  PS=1.42e-06  SA=1.9e-07  SB=9.7e-07  NRD=2.099  NRS=1.471  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M2:SRC ZN 30.5389 
R1 M7:SRC ZN 30.9166 
R2 ZN M5:SRC 31.4765 
CC44964 ZN A2 1.4821e-16
CC44962 ZN M4:GATE 4.7e-18
CC44961 ZN M5:GATE 3.83e-18
CC44960 ZN M8:GATE 4.84e-18
CC44990 ZN A1 6.208e-17
CC44992 ZN M3:GATE 3.53e-18
CC44997 ZN M2:GATE 4.44e-18
CC44972 ZN A1:1 1.532e-17
CC44978 ZN M7:GATE 7.6e-18
CC44984 ZN M6:GATE 1.018e-17
R3 M6:DRN M5:SRC 0.001 
R4 M5:SRC M7:SRC 2042.18 
CC44957 M5:SRC A2 6.8e-18
CC44956 M5:SRC M5:GATE 2.846e-17
CC44987 M5:SRC A1 1.19e-18
CC44982 M5:SRC M6:GATE 2.789e-17
R5 M7:SRC M8:DRN 0.001 
CC44959 M7:SRC A2 6.26e-18
CC44958 M7:SRC M8:GATE 2.832e-17
CC44975 M7:SRC M7:GATE 2.776e-17
R6 M2:SRC M3:DRN 0.001 
CC44988 M2:SRC A1 1.155e-17
CC44970 M2:SRC A1:1 5.852e-17
C7 ZN 0 4.694e-17
C8 M5:SRC 0 4.33e-18
C9 M7:SRC 0 4.3e-18
C10 M2:SRC 0 5.44e-18
R11 A2 M5:GATE 150.805 
R12 M5:GATE M1:GATE 469.82 
CC44983 M5:GATE M6:GATE 7.02e-18
R13 M1:GATE A2 123.522 
CC44996 M1:GATE M2:GATE 7.61e-18
CC44989 M1:GATE A1 1.073e-17
CC44971 M1:GATE A1:1 6.37e-18
R14 M4:GATE A2 118.243 
R15 A2 M8:GATE 144.361 
CC44991 A2 A1 2.937e-17
CC44985 A2 M6:GATE 8.8e-18
CC44973 A2 A1:1 3.36e-18
CC44979 A2 M7:GATE 1.093e-17
R16 M8:GATE M4:GATE 508.7 
CC44966 M8:GATE A1:1 6.42e-18
CC44974 M8:GATE M7:GATE 6.96e-18
CC44993 M4:GATE M3:GATE 1.239e-17
CC44969 M4:GATE A1:1 2.35e-18
C17 M5:GATE 0 6.728e-17
C18 M1:GATE 0 5.149e-17
C19 A2 0 3.3033e-16
C20 M8:GATE 0 5.342e-17
C21 M4:GATE 0 4.06e-17
R22 M6:GATE A1 285.883 
R23 M2:GATE A1 206.924 
R24 A1 A1:1 51.651 
R25 M6:GATE A1:1 260.68 
R26 M2:GATE A1:1 188.682 
R27 M3:GATE A1:1 94.0755 
R28 A1:1 M7:GATE 111.3 
R29 M2:GATE M6:GATE 1044.33 
C30 A1 0 1.252e-17
C31 A1:1 0 1.28e-17
C32 M7:GATE 0 4.626e-17
C33 M3:GATE 0 3.379e-17
C34 M2:GATE 0 3.469e-17
C35 M6:GATE 0 5.027e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
