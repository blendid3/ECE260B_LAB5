.SUBCKT XNR2D4 A1 A2 ZN
MMM20 M20:DRN M20:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=7.9e-14  AS=6.8e-14  PD=1.39e-06  PS=7.8e-07  SA=1.49e-07  SB=1.26e-06  NRD=0.528  NRS=0.654  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 M15:SRC M21:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.3e-14  AS=5.2e-14  PD=7.72e-07  PS=7.2e-07  SA=9.4e-07  SB=4.65e-07  NRD=4.009  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 vdd M22:GATE M22:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=8.1e-07  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 M22:SRC M23:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=1.097e-06  NRD=2.057  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 vdd M24:GATE M24:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=1.37e-06  NRD=2.099  NRS=0.427  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM25 M25:DRN M25:GATE M25:SRC vdd pch L=6e-08 W=4.5e-07  AD=6.8e-14  AS=4.5e-14  PD=1.25e-06  PS=6.5e-07  SA=4.25e-07  SB=1.48e-07  NRD=0.533  NRS=2.355  SCA=6.198  SCB=0.006  SCC=0.0002245 
MMM26 M26:DRN M26:GATE M25:SRC vdd pch L=6e-08 W=4.5e-07  AD=7.4e-14  AS=4.5e-14  PD=1.23e-06  PS=6.5e-07  SA=1.65e-07  SB=4.09e-07  NRD=0.548  NRS=2.355  SCA=6.198  SCB=0.006  SCC=0.0002245 
MMM10 M9:SRC M10:GATE vss vss nch L=6e-08 W=3.9e-07  AD=4.1e-14  AS=3.9e-14  PD=6.57e-07  PS=5.9e-07  SA=9.4e-07  SB=4.22e-07  NRD=5.786  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=7.6e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.11e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M11:SRC M12:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=1.052e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=8.46e-07  SB=4.2e-07  NRD=4.141  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.2e-14  PD=5.9e-07  PS=1.1e-06  SA=1.6e-07  SB=1.328e-06  NRD=4.183  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=5.76e-07  SB=6.8e-07  NRD=4.183  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE M14:SRC vdd pch L=6e-08 W=4.5e-07  AD=7.4e-14  AS=4.9e-14  PD=1.23e-06  PS=6.7e-07  SA=1.48e-06  SB=1.65e-07  NRD=0.548  NRS=0.313  SCA=8.144  SCB=0.009  SCC=0.0005086 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=4e-14  PD=5.9e-07  PS=6.65e-07  SA=2.85e-07  SB=9.4e-07  NRD=4.141  NRS=8.121  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 M14:SRC M15:GATE M15:SRC vdd pch L=6e-08 W=4.52e-07  AD=4.9e-14  AS=4.6e-14  PD=6.7e-07  PS=6.68e-07  SA=1.2e-06  SB=4.45e-07  NRD=0.313  NRS=0.295  SCA=8.144  SCB=0.009  SCC=0.0005086 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=3.02e-07  AD=4.8e-14  AS=2.9e-14  PD=9.1e-07  PS=4.95e-07  SA=1.65e-07  SB=1.19e-06  NRD=0.67  NRS=0.63  SCA=7.626  SCB=0.008  SCC=0.0002931 
MMM16 vdd M16:GATE M16:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.24e-06  SB=1.6e-07  NRD=0.532  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE M6:SRC vss nch L=6e-08 W=2.97e-07  AD=5.5e-14  AS=2.9e-14  PD=9.6e-07  PS=4.93e-07  SA=4.25e-07  SB=1.9e-07  NRD=1.357  NRS=3.721  SCA=7.626  SCB=0.008  SCC=0.0002931 
MMM17 M17:DRN M17:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.91e-07  SB=4.2e-07  NRD=2.057  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 M7:DRN M7:GATE M6:SRC vss nch L=6e-08 W=3.1e-07  AD=5.1e-14  AS=3.1e-14  PD=9.5e-07  PS=5.27e-07  SA=1.65e-07  SB=3.95e-07  NRD=0.643  NRS=6.111  SCA=7.393  SCB=0.008  SCC=0.0002747 
MMM18 vdd M18:GATE M18:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7.31e-07  SB=6.8e-07  NRD=2.099  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE M8:SRC vss nch L=6.1e-08 W=3.14e-07  AD=5.9e-14  AS=3.1e-14  PD=1e-06  PS=5.1e-07  SA=1.46e-06  SB=1.9e-07  NRD=1.35  NRS=5.229  SCA=8.2  SCB=0.009  SCC=0.0003833 
MMM19 M19:DRN M19:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.8e-14  PD=7.2e-07  PS=7.8e-07  SA=4.7e-07  SB=9.4e-07  NRD=2.057  NRS=0.654  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 M8:SRC M9:GATE M9:SRC vss nch L=6e-08 W=3.15e-07  AD=3.1e-14  AS=3.3e-14  PD=5.1e-07  PS=5.23e-07  SA=1.2e-06  SB=4.5e-07  NRD=5.229  NRS=0.379  SCA=8.2  SCB=0.009  SCC=0.0003833 
R0 ZN M4:DRN 15.2949 
R1 M4:DRN M3:SRC 0.001 
CC29845 M4:DRN M4:GATE 1.792e-17
CC29818 M4:DRN N_4:3 3.41e-18
CC29785 M4:DRN N_4:1 6.54e-17
CC29793 M4:DRN N_4:2 2.096e-17
CC29850 M4:DRN M3:GATE 9.9e-18
R2 M19:DRN ZN 15.3486 
R3 M17:DRN ZN 15.6708 
R4 ZN M2:DRN 15.6755 
CC29841 ZN M16:GATE 4.24e-18
CC29795 ZN N_4:2 4.69e-18
CC29857 ZN M1:GATE 5.03e-18
CC29834 ZN M18:GATE 1.258e-17
CC29828 ZN M19:GATE 4.21e-18
CC29838 ZN M17:GATE 8.67e-18
CC29819 ZN N_4:3 1.0613e-16
CC29787 ZN N_4:1 3.438e-17
CC29885 ZN M25:DRN 4.6e-18
CC29908 ZN M6:DRN 3.69e-18
CC29846 ZN M4:GATE 3.17e-18
CC29854 ZN M2:GATE 3.05e-18
CC29852 ZN M3:GATE 5.86e-18
R5 M2:DRN M1:SRC 0.001 
CC29794 M2:DRN N_4:2 4.405e-17
CC29858 M2:DRN M1:GATE 1.495e-17
CC29786 M2:DRN N_4:1 1.36e-17
CC29856 M2:DRN M2:GATE 4.164e-17
R6 M19:DRN M17:DRN 1778.96 
R7 M17:DRN M16:SRC 0.001 
CC29840 M17:DRN M16:GATE 4.701e-17
CC29837 M17:DRN M17:GATE 4.684e-17
CC29781 M17:DRN N_4:1 1.543e-17
CC29792 M17:DRN N_4:2 5.36e-18
R8 M19:DRN M18:SRC 0.001 
CC29832 M19:DRN M18:GATE 4.689e-17
CC29827 M19:DRN M19:GATE 4.708e-17
CC29805 M19:DRN N_4:3 2.87e-18
CC29780 M19:DRN N_4:1 2.055e-17
C9 M4:DRN 0 9.43e-18
C10 ZN 0 3.0384e-16
C11 M2:DRN 0 1.467e-17
C12 M17:DRN 0 2.3e-17
C13 M19:DRN 0 9.56e-18
R14 M14:DRN M15:SRC 117.159 
R15 M9:SRC M15:SRC 122.802 
R16 M15:SRC M8:DRN 127.002 
CC29702 M15:SRC M10:GATE 7.84e-18
CC29872 M15:SRC M14:SRC 8.78e-18
CC29711 M15:SRC M11:SRC 1.38e-18
CC29766 M15:SRC M14:GATE 5.51e-18
CC29753 M15:SRC M15:GATE 4.189e-17
CC29680 M15:SRC M21:GATE 3.404e-17
CC29891 M15:SRC M8:SRC 4.95e-18
CC29802 M15:SRC N_4:3 1.6e-17
CC29645 M15:SRC N_16:1 3.65e-18
CC29653 M15:SRC M8:GATE 5.95e-18
CC29669 M15:SRC N_10:2 4.789e-17
CC29651 M15:SRC M9:GATE 5.77e-18
R17 M14:DRN M8:DRN 130.657 
R18 M8:DRN M9:SRC 117.757 
CC29812 M8:DRN N_4:3 1.3072e-16
CC29758 M8:DRN M15:GATE 1.34e-18
CC29744 M8:DRN M7:GATE 2.04e-18
CC29917 M8:DRN M7:DRN 1.273e-17
CC29654 M8:DRN M8:GATE 1.107e-17
CC29648 M8:DRN N_16:1 2.366e-17
R19 M9:SRC M14:DRN 126.335 
CC29705 M9:SRC M10:GATE 9.47e-18
CC29674 M9:SRC N_10:2 1.2345e-16
CC29809 M9:SRC N_4:3 2.759e-17
CC29647 M9:SRC N_16:1 3.088e-17
CC29865 M14:DRN M26:DRN 1.309e-17
CC29670 M14:DRN N_10:2 5.08e-18
CC29768 M14:DRN M14:GATE 3.366e-17
CC29808 M14:DRN N_4:3 3.275e-17
CC29650 M14:DRN M26:GATE 1.25e-18
C20 M15:SRC 0 1.431e-17
C21 M8:DRN 0 1.948e-17
C22 M9:SRC 0 5.18e-18
C23 M14:DRN 0 1.1411e-16
R24 M13:GATE M24:GATE 1011.14 
R25 A2 M24:GATE 254.01 
R26 M24:GATE A2:1 296.35 
CC29666 M24:GATE N_10:2 7.93e-18
CC29683 M24:GATE M24:SRC 4.862e-17
R27 M12:GATE A2:1 95.3999 
R28 M22:GATE A2:1 165.597 
R29 M11:GATE A2:1 143.651 
R30 M13:GATE A2:1 237.556 
R31 A2 A2:1 59.6772 
R32 A2:1 M23:GATE 109.975 
CC29698 A2:1 M22:SRC 5.4e-18
CC29677 A2:1 N_10:2 1.501e-17
CC29714 A2:1 M11:SRC 3.753e-17
CC29709 A2:1 M10:GATE 4.5e-18
CC29667 M23:GATE N_10:2 7.52e-18
CC29694 M23:GATE M22:SRC 4.705e-17
R33 A2 M13:GATE 203.615 
CC29697 A2 M22:SRC 1.362e-17
CC29676 A2 N_10:2 8.971e-17
CC29681 A2 M21:GATE 9.8e-18
CC29701 A2 M13:SRC 3.23e-17
CC29685 A2 M24:SRC 6.65e-18
CC29671 M13:GATE N_10:2 2.116e-17
R34 M11:GATE M22:GATE 611.434 
CC29704 M11:GATE M10:GATE 4.29e-18
CC29673 M11:GATE N_10:2 3.04e-18
CC29679 M22:GATE M21:GATE 1.201e-17
CC29695 M22:GATE M22:SRC 4.698e-17
CC29668 M22:GATE N_10:2 1.406e-17
CC29712 M12:GATE M11:SRC 2.811e-17
C35 M24:GATE 0 7.826e-17
C36 A2:1 0 6.362e-17
C37 M23:GATE 0 5.881e-17
C38 A2 0 9.66e-18
C39 M13:GATE 0 5.039e-17
C40 M11:GATE 0 6.248e-17
C41 M22:GATE 0 5.089e-17
C42 M12:GATE 0 2.311e-17
R43 N_16:1 M20:DRN 192.053 
R44 M25:GATE M20:DRN 758.253 
R45 M20:DRN M5:DRN 77.0233 
CC29721 M20:DRN A1:1 4.17e-18
CC29884 M20:DRN M25:DRN 3.79e-18
CC29862 M20:DRN M26:DRN 1.01e-18
CC29749 M20:DRN M5:GATE 5.74e-18
CC29754 M20:DRN M15:GATE 5.33e-18
CC29902 M20:DRN M6:DRN 4.92e-18
CC29767 M20:DRN M14:GATE 1.482e-17
CC29732 M20:DRN M20:GATE 2.91e-18
CC29737 M20:DRN A1 1.0331e-16
CC29742 M20:DRN M7:GATE 3.036e-17
CC29804 M20:DRN N_4:3 6.94e-18
R46 N_16:1 M5:DRN 194.471 
R47 M5:DRN M25:GATE 767.806 
CC29727 M5:DRN A1:1 2.05e-18
CC29750 M5:DRN M5:GATE 7.58e-18
CC29907 M5:DRN M6:DRN 8.62e-18
CC29759 M5:DRN M15:GATE 3.09e-18
CC29739 M5:DRN A1 2.257e-17
CC29662 M5:DRN N_10:1 7.74e-17
CC29746 M5:DRN M7:GATE 1.548e-17
CC29817 M5:DRN N_4:3 6.751e-17
R48 M25:GATE N_16:1 190.392 
CC29688 M25:GATE M25:SRC 5.27e-18
CC29882 M25:GATE M25:DRN 2.963e-17
CC29798 M25:GATE N_4:3 9.94e-18
CC29656 M25:GATE N_10:1 1.142e-17
R49 M9:GATE N_16:1 235.025 
R50 M8:GATE N_16:1 130.858 
R51 N_16:1 M26:GATE 108.651 
CC29692 N_16:1 M25:SRC 6.197e-17
CC29868 N_16:1 M26:DRN 3e-18
CC29822 N_16:1 N_4:3 1.3452e-16
CC29747 N_16:1 M7:GATE 9.39e-18
CC29910 N_16:1 M6:DRN 1.28e-18
CC29771 N_16:1 M14:GATE 2.85e-18
CC29761 N_16:1 M15:GATE 1.85e-18
CC29899 N_16:1 M8:SRC 3.942e-17
CC29920 N_16:1 M7:DRN 3.32e-18
CC29888 N_16:1 M25:DRN 3.32e-18
CC29878 N_16:1 M14:SRC 2.54e-18
CC29717 N_16:1 M6:SRC 2.14e-18
CC29710 N_16:1 M10:GATE 3.8e-18
CC29860 M26:GATE M26:DRN 2.909e-17
CC29687 M26:GATE M25:SRC 4.01e-17
CC29763 M26:GATE M14:GATE 1.62e-18
CC29664 M26:GATE N_10:2 4.58e-18
CC29797 M26:GATE N_4:3 3.11e-18
CC29655 M26:GATE N_10:1 2.1e-18
R52 M8:GATE M9:GATE 319.997 
CC29757 M8:GATE M15:GATE 3.257e-17
CC29811 M8:GATE N_4:3 5.366e-17
CC29724 M9:GATE A1:1 3.95e-18
CC29896 M9:GATE M8:SRC 3.047e-17
CC29661 M9:GATE N_10:1 3.816e-17
CC29706 M9:GATE M10:GATE 4.14e-18
CC29810 M9:GATE N_4:3 1.89e-18
C53 M20:DRN 0 2.554e-17
C54 M5:DRN 0 1.424e-17
C55 M25:GATE 0 3.588e-17
C56 N_16:1 0 8.55e-18
C57 M26:GATE 0 2.432e-17
C58 M8:GATE 0 2.287e-17
C59 M9:GATE 0 2.396e-17
R60 M22:SRC N_10:1 94.5924 
R61 M24:SRC N_10:1 118.586 
R62 N_10:2 N_10:1 3.67552 
R63 M6:SRC N_10:1 31.5206 
R64 N_10:1 M25:SRC 15.1445 
CC29772 N_10:1 M14:GATE 6.21e-18
CC29823 N_10:1 N_4:3 8.503e-17
CC29879 N_10:1 M14:SRC 1.341e-17
CC29889 N_10:1 M25:DRN 1.12e-18
CC29869 N_10:1 M26:DRN 1.769e-17
CC29729 N_10:1 A1:1 5.49e-18
CC29748 N_10:1 M7:GATE 1.02e-17
CC29740 N_10:1 A1 1.17e-18
R65 M25:SRC M6:SRC 3192.69 
CC29796 M25:SRC N_4:3 2.35e-18
CC29814 M6:SRC N_4:3 4.7e-18
CC29726 M6:SRC A1:1 5.499e-17
CC29745 M6:SRC M7:GATE 2.037e-17
R66 M10:GATE M21:GATE 538.048 
R67 M21:GATE N_10:2 147.759 
CC29801 M21:GATE N_4:3 1.95e-18
CC29752 M21:GATE M15:GATE 6.82e-18
R68 M22:SRC N_10:2 18.7587 
R69 M11:SRC N_10:2 31.0107 
R70 M13:SRC N_10:2 31.8549 
R71 M10:GATE N_10:2 121.901 
R72 N_10:2 M24:SRC 18.7257 
CC29867 N_10:2 M26:DRN 3.04e-18
CC29821 N_10:2 N_4:3 1.52e-18
CC29877 N_10:2 M14:SRC 2.57e-18
CC29760 N_10:2 M15:GATE 1.029e-17
CC29799 M24:SRC N_4:3 1.034e-17
R73 M13:SRC M11:SRC 1866.06 
CC29800 M22:SRC N_4:3 1.65e-18
C74 N_10:1 0 9e-17
C75 M25:SRC 0 5.48e-18
C76 M6:SRC 0 6.76e-18
C77 M21:GATE 0 3.649e-17
C78 N_10:2 0 3.2446e-16
C79 M24:SRC 0 2.083e-17
C80 M10:GATE 0 3.345e-17
C81 M13:SRC 0 1.622e-17
C82 M11:SRC 0 7.9e-18
C83 M22:SRC 0 1.969e-17
R84 M5:GATE A1 143.889 
R85 M20:GATE A1 170.009 
R86 A1 A1:1 251.1 
CC29886 A1 M25:DRN 2.84e-18
CC29788 A1 N_4:1 2.13e-18
CC29820 A1 N_4:3 4.38e-17
CC29829 A1 M19:GATE 5.76e-18
R87 M6:GATE A1:1 67.5751 
R88 M14:GATE A1:1 883.513 
R89 M7:GATE A1:1 158.338 
R90 M15:GATE A1:1 1589 
R91 M5:GATE A1:1 427.502 
R92 A1:1 M20:GATE 1222.64 
CC29912 A1:1 M6:DRN 1.098e-17
CC29922 A1:1 M7:DRN 3.96e-17
CC29870 A1:1 M26:DRN 1.65e-18
CC29790 A1:1 N_4:1 1.44e-18
CC29824 A1:1 N_4:3 7.77e-18
R93 M20:GATE M5:GATE 700.614 
CC29883 M20:GATE M25:DRN 1.73e-18
CC29803 M20:GATE N_4:3 8.81e-18
CC29778 M20:GATE N_4:1 1.72e-18
CC29906 M5:GATE M6:DRN 2.17e-18
CC29844 M5:GATE M4:GATE 4.34e-18
CC29816 M5:GATE N_4:3 5.62e-18
CC29783 M5:GATE N_4:1 1.212e-17
R94 M14:GATE M15:GATE 310.183 
R95 M15:GATE M7:GATE 1619.56 
CC29892 M15:GATE M8:SRC 1e-18
CC29874 M15:GATE M14:SRC 3.797e-17
CC29806 M15:GATE N_4:3 1.238e-17
R96 M7:GATE M14:GATE 900.505 
CC29813 M7:GATE N_4:3 5.27e-18
CC29893 M14:GATE M8:SRC 9.47e-18
CC29875 M14:GATE M14:SRC 2.893e-17
CC29864 M14:GATE M26:DRN 4.87e-18
CC29915 M14:GATE M7:DRN 4.27e-18
CC29807 M14:GATE N_4:3 4.63e-18
CC29782 M14:GATE N_4:1 1.61e-18
CC29905 M6:GATE M6:DRN 2.278e-17
CC29815 M6:GATE N_4:3 2.5e-18
C97 A1 0 2.97e-18
C98 A1:1 0 7.26e-18
C99 M20:GATE 0 4.3e-17
C100 M5:GATE 0 2.636e-17
C101 M15:GATE 0 2.629e-17
C102 M7:GATE 0 3.275e-17
C103 M14:GATE 0 3.585e-17
C104 M6:GATE 0 2.211e-17
R105 M17:GATE N_4:2 106 
R106 M2:GATE N_4:2 99.3746 
R107 M1:GATE N_4:2 146.49 
R108 M16:GATE N_4:2 156.256 
R109 M3:GATE N_4:2 254.147 
R110 M18:GATE N_4:2 271.09 
R111 N_4:2 N_4:1 57.4072 
R112 M19:GATE N_4:1 106 
R113 M6:DRN N_4:1 720.66 
R114 M4:GATE N_4:1 90.365 
R115 M3:GATE N_4:1 234.598 
R116 M18:GATE N_4:1 250.238 
R117 N_4:3 N_4:1 27.778 
R118 N_4:1 M25:DRN 301.856 
R119 M6:DRN M25:DRN 1034.27 
R120 M25:DRN N_4:3 39.8663 
R121 M7:DRN N_4:3 29.9999 
R122 M6:DRN N_4:3 33.5244 
R123 M8:SRC N_4:3 32.3801 
R124 M14:SRC N_4:3 34.3734 
R125 N_4:3 M26:DRN 35.2456 
R126 M8:SRC M26:DRN 1270.97 
R127 M26:DRN M14:SRC 589.767 
R128 M14:SRC M8:SRC 1239.51 
R129 M18:GATE M3:GATE 1107.81 
R130 M16:GATE M1:GATE 638.548 
C131 M17:GATE 0 4.802e-17
C132 N_4:2 0 3.991e-17
C133 N_4:1 0 7.174e-17
C134 M25:DRN 0 5.061e-17
C135 N_4:3 0 1.073e-16
C136 M26:DRN 0 7.54e-18
C137 M14:SRC 0 7.85e-18
C138 M8:SRC 0 7.82e-18
C139 M18:GATE 0 5.507e-17
C140 M3:GATE 0 5.766e-17
C141 M16:GATE 0 8.405e-17
C142 M1:GATE 0 6.192e-17
C143 M4:GATE 0 2.763e-17
C144 M2:GATE 0 2.063e-17
C145 M6:DRN 0 3.537e-17
C146 M19:GATE 0 4.761e-17
C147 M7:DRN 0 9.58e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
