.SUBCKT BUFFD16 I Z
MMM20 M19:SRC M20:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.35e-07  SB=5.145e-06  NRD=4.183  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM21 M21:DRN M21:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.8e-14  AS=3.9e-14  PD=1.13e-06  PS=5.9e-07  SA=1.75e-07  SB=5.405e-06  NRD=0.592  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM22 vdd M22:GATE M22:SRC vdd pch L=6e-08 W=5.2e-07  AD=1.07e-13  AS=5.2e-14  PD=1.45e-06  PS=7.2e-07  SA=5.375e-06  SB=2.05e-07  NRD=0.488  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 M23:DRN M23:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=5.115e-06  SB=4.65e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 vdd M24:GATE M24:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.855e-06  SB=7.25e-07  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM25 M25:DRN M25:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.595e-06  SB=9.85e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM26 vdd M26:GATE M26:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.335e-06  SB=1.245e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM27 M27:DRN M27:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.075e-06  SB=1.505e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM28 vdd M28:GATE M28:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.815e-06  SB=1.765e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM29 M29:DRN M29:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.555e-06  SB=2.025e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM40 vdd M40:GATE M40:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.95e-07  SB=4.885e-06  NRD=2.534  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM41 M40:SRC M41:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.35e-07  SB=5.145e-06  NRD=2.099  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM42 M42:DRN M42:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=9.1e-14  AS=5.2e-14  PD=1.39e-06  PS=7.2e-07  SA=1.75e-07  SB=5.405e-06  NRD=0.541  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.035e-06  SB=2.545e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.775e-06  SB=2.805e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=8e-14  AS=3.9e-14  PD=1.19e-06  PS=5.9e-07  SA=5.375e-06  SB=2.05e-07  NRD=0.566  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.515e-06  SB=3.065e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=5.115e-06  SB=4.65e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.255e-06  SB=3.325e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.855e-06  SB=7.25e-07  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.995e-06  SB=3.585e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.595e-06  SB=9.85e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vss M15:GATE M15:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.735e-06  SB=3.845e-06  NRD=4.537  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.335e-06  SB=1.245e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.475e-06  SB=4.105e-06  NRD=4.183  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.075e-06  SB=1.505e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 vss M17:GATE M17:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.215e-06  SB=4.365e-06  NRD=4.537  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.815e-06  SB=1.765e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M17:SRC M18:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.55e-07  SB=4.625e-06  NRD=4.183  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.555e-06  SB=2.025e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vss M19:GATE M19:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.95e-07  SB=4.885e-06  NRD=4.537  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.295e-06  SB=2.285e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM30 vdd M30:GATE M30:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.295e-06  SB=2.285e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM31 M31:DRN M31:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.035e-06  SB=2.545e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM32 vdd M32:GATE M32:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.775e-06  SB=2.805e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM33 M33:DRN M33:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.515e-06  SB=3.065e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM34 vdd M34:GATE M34:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.255e-06  SB=3.325e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM35 M35:DRN M35:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.995e-06  SB=3.585e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM36 vdd M36:GATE M36:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.735e-06  SB=3.845e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM37 M37:DRN M37:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.475e-06  SB=4.105e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM38 vdd M38:GATE M38:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.215e-06  SB=4.365e-06  NRD=2.534  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM39 M38:SRC M39:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.55e-07  SB=4.625e-06  NRD=2.099  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M27:DRN Z:3 41.6887 
R1 Z:1 Z:3 0.50175 
R2 M29:DRN Z:3 20.6283 
R3 M31:DRN Z:3 14.9999 
R4 M34:SRC Z:3 16.0439 
R5 M33:DRN Z:3 15.6689 
R6 M37:DRN Z:3 16.2369 
R7 Z:3 Z 0.104 
CC30018 Z:3 M31:GATE 1.794e-17
CC29991 Z:3 N_10:3 1.0465e-16
CC30012 Z:3 M32:GATE 1.685e-17
CC30009 Z:3 M40:SRC 6.95e-18
CC30001 Z:3 N_10:6 1.0659e-16
CC30112 Z:3 N_10:15 4.592e-17
CC30171 Z:3 M38:SRC 4.12e-18
CC30039 Z:3 M26:GATE 1.82e-17
CC30044 Z:3 M25:GATE 1.782e-17
CC30048 Z:3 M24:GATE 1.82e-17
CC30053 Z:3 M23:GATE 1.704e-17
CC30022 Z:3 M30:GATE 1.461e-17
CC30026 Z:3 M29:GATE 1.657e-17
CC30030 Z:3 M28:GATE 1.767e-17
CC30035 Z:3 M27:GATE 1.743e-17
CC30057 Z:3 M22:GATE 4.83e-18
CC30207 Z:3 M33:GATE 1.885e-17
CC30202 Z:3 M34:GATE 1.659e-17
CC30197 Z:3 M35:GATE 1.839e-17
CC30192 Z:3 M36:GATE 1.565e-17
CC30187 Z:3 M37:GATE 4.58e-18
CC30182 Z:3 M42:DRN 6.73e-18
R8 Z Z:2 0.09776 
R9 M6:DRN Z:2 15.6919 
R10 M8:DRN Z:2 15.0384 
R11 M10:DRN Z:2 14.9999 
R12 M4:DRN Z:2 16.0794 
R13 M13:SRC Z:2 15.4941 
R14 M15:SRC Z:2 31.1808 
R15 M12:DRN Z:2 15.3585 
R16 Z:2 M2:DRN 16.2792 
CC30019 Z:2 M31:GATE 3.91e-18
CC29992 Z:2 N_10:3 1.5187e-16
CC29961 Z:2 N_10:1 3.36e-18
CC29965 Z:2 N_10:2 5.65e-18
CC30002 Z:2 N_10:6 1.4705e-16
CC30013 Z:2 M32:GATE 1.78e-18
CC30126 Z:2 M10:GATE 1.16e-17
CC30121 Z:2 M11:GATE 1.23e-17
CC30120 Z:2 N_10:16 2.11e-18
CC30113 Z:2 N_10:15 9.647e-17
CC30090 Z:2 N_10:14 2.39e-18
CC30145 Z:2 M3:GATE 1.242e-17
CC30148 Z:2 M2:GATE 1.224e-17
CC30152 Z:2 M1:GATE 3.61e-18
CC30153 Z:2 M14:GATE 1.49e-17
CC30156 Z:2 M15:GATE 1.217e-17
CC30165 Z:2 M16:GATE 4.87e-18
CC30129 Z:2 M9:GATE 1.123e-17
CC30132 Z:2 M8:GATE 1.603e-17
CC30135 Z:2 M7:GATE 1.168e-17
CC30136 Z:2 M6:GATE 1.246e-17
CC30141 Z:2 M5:GATE 1.246e-17
CC30142 Z:2 M4:GATE 1.246e-17
CC30023 Z:2 M30:GATE 6.8e-18
CC30027 Z:2 M29:GATE 2.53e-18
CC30031 Z:2 M28:GATE 1.91e-18
CC30071 Z:2 N_10:9 1.85e-18
CC30075 Z:2 N_10:10 2.93e-18
CC30076 Z:2 N_10:11 2.94e-18
CC30082 Z:2 N_10:12 3.08e-18
CC30086 Z:2 N_10:13 2.93e-18
CC30062 Z:2 N_10:7 3.02e-18
CC30067 Z:2 N_10:8 1.43e-18
CC30221 Z:2 M13:GATE 1.211e-17
CC30224 Z:2 M12:GATE 4.65e-18
CC30177 Z:2 M17:SRC 2.77e-18
R17 M6:DRN M2:DRN 1037.57 
R18 M4:DRN M2:DRN 575.056 
R19 M2:DRN M1:SRC 0.001 
CC30000 M2:DRN N_10:6 1.697e-17
CC30107 M2:DRN N_10:15 1.386e-17
CC30150 M2:DRN M2:GATE 5.45e-18
CC30151 M2:DRN M1:GATE 5.32e-18
CC30084 M2:DRN N_10:13 6.897e-17
R20 M12:DRN M11:SRC 0.001 
CC29985 M12:DRN N_10:3 1.36e-18
CC30122 M12:DRN M11:GATE 1.127e-17
CC30102 M12:DRN N_10:15 4.761e-17
CC30068 M12:DRN N_10:9 3.689e-17
CC30225 M12:DRN M12:GATE 1.431e-17
R21 M16:DRN M15:SRC 0.001 
R22 M15:SRC M13:SRC 1416.81 
CC29968 M15:SRC N_10:3 9.98e-18
CC29983 M15:SRC N_10:3 2.29e-18
CC30114 M15:SRC N_10:16 4.004e-17
CC30100 M15:SRC N_10:15 1.036e-17
CC30161 M15:SRC M16:GATE 6.15e-18
R23 M13:SRC M14:DRN 0.001 
CC29984 M13:SRC N_10:3 1.34e-18
CC30088 M13:SRC N_10:14 4.127e-17
CC30101 M13:SRC N_10:15 1.442e-17
CC30155 M13:SRC M14:GATE 6.24e-18
CC30064 M13:SRC N_10:8 3.954e-17
CC30223 M13:SRC M13:GATE 8.29e-18
R24 M36:SRC M37:DRN 0.001 
R25 M34:SRC M37:DRN 593.061 
R26 M37:DRN M33:DRN 1071.03 
CC29975 M37:DRN N_10:3 2.45e-18
CC30092 M37:DRN N_10:15 1.234e-17
CC30189 M37:DRN M36:GATE 4.554e-17
CC30185 M37:DRN M37:GATE 4.607e-17
R27 M32:SRC M33:DRN 0.001 
R28 M33:DRN M34:SRC 1058.29 
CC30010 M33:DRN M32:GATE 4.555e-17
CC29977 M33:DRN N_10:3 1.4e-18
CC30094 M33:DRN N_10:15 1.163e-17
CC30206 M33:DRN M33:GATE 4.603e-17
R29 M34:SRC M35:DRN 0.001 
CC29976 M34:SRC N_10:3 1.4e-18
CC30093 M34:SRC N_10:15 1.163e-17
CC30200 M34:SRC M34:GATE 4.556e-17
CC30195 M34:SRC M35:GATE 4.616e-17
R30 M6:DRN M4:DRN 1024.84 
R31 M4:DRN M3:SRC 0.001 
CC29999 M4:DRN N_10:6 1.07e-18
CC30106 M4:DRN N_10:15 1.409e-17
CC30144 M4:DRN M4:GATE 7.82e-18
CC30146 M4:DRN M3:GATE 7.5e-18
CC30078 M4:DRN N_10:11 4.045e-17
CC30079 M4:DRN N_10:12 4.108e-17
R32 M31:DRN M30:SRC 0.001 
CC30015 M31:DRN M31:GATE 4.521e-17
CC30095 M31:DRN N_10:15 1.158e-17
CC30020 M31:DRN M30:GATE 4.49e-17
R33 M28:SRC M29:DRN 0.001 
R34 M29:DRN Z:1 56.307 
CC30096 M29:DRN N_10:15 1.172e-17
CC30025 M29:DRN M29:GATE 4.543e-17
CC30028 M29:DRN M28:GATE 4.547e-17
R35 M23:DRN Z:1 15.1806 
R36 M25:DRN Z:1 14.9999 
R37 Z:1 M27:DRN 23.8319 
R38 M27:DRN M26:SRC 0.001 
CC29994 M27:DRN N_10:6 1.4e-18
CC30097 M27:DRN N_10:15 1.163e-17
CC30037 M27:DRN M26:GATE 4.593e-17
CC30034 M27:DRN M27:GATE 4.567e-17
R39 M25:DRN M24:SRC 0.001 
CC29995 M25:DRN N_10:6 1.4e-18
CC30098 M25:DRN N_10:15 1.163e-17
CC30043 M25:DRN M25:GATE 4.567e-17
CC30046 M25:DRN M24:GATE 4.594e-17
R40 M10:DRN M9:SRC 0.001 
CC29963 M10:DRN N_10:2 5.409e-17
CC30125 M10:DRN M10:GATE 1.481e-17
CC30103 M10:DRN N_10:15 1.403e-17
CC30127 M10:DRN M9:GATE 9.95e-18
CC30069 M10:DRN N_10:9 1.599e-17
R41 M23:DRN M22:SRC 0.001 
CC29996 M23:DRN N_10:6 1.34e-18
CC30099 M23:DRN N_10:15 1.146e-17
CC30052 M23:DRN M23:GATE 4.496e-17
CC30056 M23:DRN M22:GATE 4.607e-17
R42 M8:DRN M7:SRC 0.001 
CC29958 M8:DRN N_10:1 5.766e-17
CC29964 M8:DRN N_10:2 1.762e-17
CC30104 M8:DRN N_10:15 1.42e-17
CC30131 M8:DRN M8:GATE 1.067e-17
CC30133 M8:DRN M7:GATE 9.83e-18
R43 M6:DRN M5:SRC 0.001 
CC29998 M6:DRN N_10:6 1.07e-18
CC30105 M6:DRN N_10:15 1.409e-17
CC30138 M6:DRN M6:GATE 5.85e-18
CC30139 M6:DRN M5:GATE 5.85e-18
CC30072 M6:DRN N_10:10 4.136e-17
CC30059 M6:DRN N_10:7 4.205e-17
C44 Z:3 0 3.7541e-16
C45 Z 0 5.6e-19
C46 Z:2 0 3.6968e-16
C47 M2:DRN 0 7.65e-18
C48 M12:DRN 0 1.439e-17
C49 M15:SRC 0 3.7e-18
C50 M13:SRC 0 5.26e-18
C51 M37:DRN 0 8.3e-18
C52 M33:DRN 0 2.093e-17
C53 M34:SRC 0 7.87e-18
C54 M4:DRN 0 2.06e-18
C55 M31:DRN 0 8.07e-18
C56 M29:DRN 0 6.75e-18
C57 M27:DRN 0 6.89e-18
C58 M25:DRN 0 7.09e-18
C59 M10:DRN 0 4.61e-18
C60 M23:DRN 0 1.146e-17
C61 M8:DRN 0 3.88e-18
C62 M6:DRN 0 4.18e-18
R63 I:2 I 56.1586 
R64 M38:GATE I 438.303 
R65 M17:GATE I 370.469 
R66 I I:3 22.8979 
CC30117 I N_10:16 2.76e-18
CC30162 I M16:GATE 1.82e-18
CC30174 I M17:SRC 1.518e-17
CC29987 I N_10:3 8.426e-17
R67 M39:GATE I:3 111.3 
R68 M18:GATE I:3 94.0755 
R69 I:2 I:3 31.0374 
R70 M38:GATE I:3 239.804 
R71 I:3 M17:GATE 202.693 
CC29990 I:3 N_10:3 1.75e-18
CC30176 I:3 M17:SRC 4.031e-17
R72 M17:GATE M38:GATE 728.434 
CC30160 M17:GATE M16:GATE 3.64e-18
CC29967 M17:GATE N_10:3 7.47e-18
CC29982 M17:GATE N_10:3 1.272e-17
CC30168 M38:GATE M38:SRC 2.762e-17
CC29974 M38:GATE N_10:3 1.294e-17
CC30184 M38:GATE M37:GATE 1.327e-17
R73 M21:GATE I:1 94.0755 
R74 M20:GATE I:1 233.022 
R75 M41:GATE I:1 275.689 
R76 M42:GATE I:1 111.3 
R77 I:1 I:2 60.2341 
CC30110 I:1 N_10:15 5.41e-18
CC30170 I:1 M38:SRC 8.9e-18
CC30008 I:1 M40:SRC 9.29e-18
CC29988 I:1 N_10:3 3.178e-17
CC30210 I:1 M21:DRN 2.644e-17
CC30217 I:1 M19:SRC 2.425e-17
CC30175 I:1 M17:SRC 1.118e-17
R78 M20:GATE I:2 233.022 
R79 M41:GATE I:2 275.689 
R80 M40:GATE I:2 111.3 
R81 I:2 M19:GATE 94.0755 
CC29989 I:2 N_10:3 1.49e-18
CC30218 I:2 M19:SRC 3.682e-17
CC29980 M19:GATE N_10:3 1.181e-17
CC30173 M18:GATE M17:SRC 1.04e-18
CC29981 M18:GATE N_10:3 1.139e-17
CC30005 M40:GATE M40:SRC 2.73e-17
CC29972 M40:GATE N_10:3 1.315e-17
CC30167 M39:GATE M38:SRC 2.766e-17
CC29973 M39:GATE N_10:3 1.142e-17
CC29970 M42:GATE N_10:3 1.299e-17
CC30178 M42:GATE M42:DRN 2.758e-17
R82 M41:GATE M20:GATE 1066.52 
CC30004 M41:GATE M40:SRC 2.73e-17
CC29971 M41:GATE N_10:3 1.481e-17
CC30212 M41:GATE M19:SRC 1.5e-18
CC29979 M20:GATE N_10:3 1.252e-17
CC30214 M20:GATE M19:SRC 3.64e-18
CC29978 M21:GATE N_10:3 1.177e-17
CC30209 M21:GATE M21:DRN 1.37e-18
C83 I 0 6.81e-18
C84 I:3 0 4.75e-18
C85 M17:GATE 0 2.582e-17
C86 M38:GATE 0 4.139e-17
C87 I:1 0 3.625e-17
C88 I:2 0 3.48e-18
C89 M19:GATE 0 3.157e-17
C90 M18:GATE 0 2.59e-17
C91 M40:GATE 0 4.221e-17
C92 M39:GATE 0 3.64e-17
C93 M42:GATE 0 3.984e-17
C94 M41:GATE 0 3.643e-17
C95 M20:GATE 0 2.636e-17
C96 M21:GATE 0 3.635e-17
R97 M30:GATE N_10:2 106 
R98 M9:GATE N_10:2 99.3746 
R99 M8:GATE N_10:2 245.865 
R100 M29:GATE N_10:2 262.256 
R101 M10:GATE N_10:2 231.204 
R102 M31:GATE N_10:2 246.616 
R103 N_10:1 N_10:2 60.1649 
R104 N_10:2 N_10:9 66.3689 
R105 M11:GATE N_10:9 85.86 
R106 N_10:15 N_10:9 22.6646 
R107 N_10:3 N_10:9 22.7252 
R108 M10:GATE N_10:9 271.218 
R109 M31:GATE N_10:9 289.302 
R110 N_10:9 M32:GATE 106 
R111 N_10:7 N_10:1 35.6744 
R112 M7:GATE N_10:1 99.3746 
R113 M8:GATE N_10:1 245.865 
R114 M29:GATE N_10:1 262.256 
R115 M28:GATE N_10:1 106 
R116 N_10:1 N_10:6 45.926 
R117 N_10:10 N_10:6 22.6603 
R118 N_10:11 N_10:6 22 
R119 M22:GATE N_10:6 267.533 
R120 M1:GATE N_10:6 216.702 
R121 N_10:12 N_10:6 22.7118 
R122 N_10:7 N_10:6 18.2745 
R123 N_10:6 N_10:13 16.4604 
R124 M2:GATE N_10:13 88.1128 
R125 M22:GATE N_10:13 258.574 
R126 M1:GATE N_10:13 209.445 
R127 N_10:12 N_10:13 22.6689 
R128 N_10:13 M23:GATE 106 
R129 M31:GATE M10:GATE 1007.81 
R130 M29:GATE M8:GATE 1071.73 
R131 M16:GATE N_10:3 210.716 
R132 M37:GATE N_10:3 226.976 
R133 N_10:16 N_10:3 15.9377 
R134 N_10:14 N_10:3 22.2409 
R135 N_10:8 N_10:3 22 
R136 N_10:15 N_10:3 22.4793 
R137 M38:SRC N_10:3 31.7084 
R138 M42:DRN N_10:3 33.1278 
R139 M40:SRC N_10:3 32.6431 
R140 M19:SRC N_10:3 32.2663 
R141 M21:DRN N_10:3 32.7461 
R142 N_10:3 M17:SRC 31.3418 
R143 M19:SRC M17:SRC 2112.7 
R144 M17:SRC M21:DRN 2144.09 
R145 M21:DRN M19:SRC 1078.6 
R146 M38:SRC M40:SRC 1678.81 
R147 M40:SRC M42:DRN 957.931 
R148 M42:DRN M38:SRC 1703.74 
R149 M33:GATE N_10:15 83.475 
R150 N_10:8 N_10:15 22.9146 
R151 N_10:15 M12:GATE 88.1128 
R152 M34:GATE N_10:8 98.4912 
R153 M13:GATE N_10:8 91.8666 
R154 N_10:8 N_10:14 21.5119 
R155 N_10:16 N_10:14 22.8293 
R156 M35:GATE N_10:14 98.4912 
R157 N_10:14 M14:GATE 91.8666 
R158 M36:GATE N_10:16 94.7372 
R159 M15:GATE N_10:16 88.1128 
R160 M16:GATE N_10:16 219.478 
R161 N_10:16 M37:GATE 236.414 
R162 M37:GATE M16:GATE 885.822 
R163 M6:GATE N_10:7 85.86 
R164 N_10:10 N_10:7 22.6035 
R165 N_10:7 M27:GATE 106 
R166 N_10:11 N_10:12 21.5119 
R167 M3:GATE N_10:12 91.8666 
R168 N_10:12 M24:GATE 106 
R169 M1:GATE M22:GATE 989.753 
R170 M4:GATE N_10:11 91.8666 
R171 N_10:10 N_10:11 22.9146 
R172 N_10:11 M25:GATE 106 
R173 M5:GATE N_10:10 88.1128 
R174 N_10:10 M26:GATE 106 
C175 M30:GATE 0 3.393e-17
C176 N_10:2 0 3.55e-18
C177 N_10:9 0 2.07e-18
C178 M32:GATE 0 1.61e-17
C179 N_10:1 0 3.81e-18
C180 N_10:6 0 6.951e-17
C181 N_10:13 0 5.15e-18
C182 M23:GATE 0 4.173e-17
C183 M28:GATE 0 2.629e-17
C184 M31:GATE 0 3.015e-17
C185 M10:GATE 0 2.385e-17
C186 M29:GATE 0 3.233e-17
C187 M8:GATE 0 2.499e-17
C188 N_10:3 0 1.8158e-16
C189 M17:SRC 0 4.56e-18
C190 M21:DRN 0 1.191e-17
C191 M19:SRC 0 6.43e-18
C192 M40:SRC 0 2.74e-18
C193 M42:DRN 0 1.638e-17
C194 M38:SRC 0 2.74e-18
C195 M33:GATE 0 3.747e-17
C196 N_10:15 0 1.2605e-16
C197 M12:GATE 0 2.913e-17
C198 M34:GATE 0 3.291e-17
C199 N_10:8 0 3.13e-18
C200 N_10:14 0 3.24e-18
C201 M14:GATE 0 2.149e-17
C202 M35:GATE 0 3.204e-17
C203 M36:GATE 0 3.513e-17
C204 N_10:16 0 2.59e-18
C205 M37:GATE 0 4.059e-17
C206 M16:GATE 0 2.895e-17
C207 M7:GATE 0 2.231e-17
C208 N_10:7 0 1.208e-17
C209 M27:GATE 0 3.179e-17
C210 M9:GATE 0 3.013e-17
C211 N_10:12 0 2.54e-18
C212 M24:GATE 0 3.03e-17
C213 M1:GATE 0 6.112e-17
C214 M22:GATE 0 8.259e-17
C215 M2:GATE 0 3.926e-17
C216 M3:GATE 0 2.519e-17
C217 M4:GATE 0 2.18e-17
C218 N_10:11 0 3.39e-18
C219 M25:GATE 0 2.644e-17
C220 M5:GATE 0 2.541e-17
C221 N_10:10 0 6.17e-18
C222 M26:GATE 0 2.961e-17
C223 M6:GATE 0 2.698e-17
C224 M11:GATE 0 1.481e-17
C225 M13:GATE 0 2.438e-17
C226 M15:GATE 0 2.734e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
