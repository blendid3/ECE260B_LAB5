.SUBCKT NR2D8 A1 A2 ZN
MMM20 M20:DRN M20:GATE M20:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.26e-06  SB=9.4e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 M20:SRC M21:GATE M21:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3e-06  SB=1.2e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE M22:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.74e-06  SB=1.46e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 M22:SRC M23:GATE M23:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.48e-06  SB=1.72e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 M24:DRN M24:GATE M24:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.22e-06  SB=1.98e-06  NRD=2.099  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM25 M24:SRC M25:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.98e-06  SB=2.22e-06  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM26 vdd M26:GATE M26:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=1.72e-06  SB=2.48e-06  NRD=6.61  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM27 M26:SRC M27:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.46e-06  SB=2.74e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM28 vdd M28:GATE M28:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.2e-06  SB=3e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM29 M28:SRC M29:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.4e-07  SB=3.26e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=1.7e-06  SB=2.5e-06  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=1.46e-06  SB=2.74e-06  NRD=7.648  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=4.04e-06  SB=1.6e-07  NRD=0.462  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.2e-06  SB=3e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.78e-06  SB=4.2e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.4e-07  SB=3.26e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.52e-06  SB=6.8e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=3.52e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.26e-06  SB=9.4e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vss M15:GATE M15:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=3.78e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3e-06  SB=1.2e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 vss M16:GATE M16:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.6e-07  SB=4.065e-06  NRD=0.567  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.74e-06  SB=1.46e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 M17:DRN M17:GATE M17:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=4.04e-06  SB=1.6e-07  NRD=0.427  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.48e-06  SB=1.72e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M18:DRN M18:GATE M18:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.78e-06  SB=4.2e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.24e-06  SB=1.985e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 M18:SRC M19:GATE M19:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.52e-06  SB=6.8e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.98e-06  SB=2.245e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM30 vdd M30:GATE M30:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=3.52e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM31 M30:SRC M31:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=3.78e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM32 vdd M32:GATE M32:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=4.04e-06  NRD=2.099  NRS=0.427  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M29:GATE A2:3 111.3 
R1 M13:GATE A2:3 83.3024 
R2 A2 A2:3 22.159 
R3 A2:4 A2:3 23.85 
R4 A2:3 A2:2 23.7579 
CC47924 A2:3 ZN:3 3.83e-18
CC47939 A2:3 M13:SRC 2.874e-17
CC48132 A2:3 M28:SRC 3.9e-18
R5 M30:GATE A2:2 111.3 
R6 M15:GATE A2:2 220.731 
R7 M14:GATE A2:2 84.4211 
R8 A2 A2:2 22.3605 
R9 A2:1 A2:2 57.0569 
R10 A2:2 M31:GATE 261.147 
CC47933 A2:2 M15:SRC 1.619e-17
CC47938 A2:2 M13:SRC 2.06e-17
CC47923 A2:2 ZN:3 1.15e-18
CC48120 A2:2 M30:SRC 8.19e-18
R11 M15:GATE M31:GATE 1108.31 
R12 M31:GATE A2:1 286.489 
CC47911 M31:GATE ZN:3 1.01e-18
CC48112 M31:GATE M30:SRC 2.592e-17
CC48136 M31:GATE N_9:3 6.97e-18
R13 M32:GATE A2:1 111.3 
R14 M15:GATE A2:1 242.151 
R15 A2:1 M16:GATE 94.0755 
CC47931 A2:1 M15:SRC 1.831e-17
CC48158 A2:1 N_9:3 1.66e-18
CC47929 M16:GATE M15:SRC 2.459e-17
CC47912 M16:GATE ZN:3 1.8e-18
R16 M12:GATE A2:4 82.3623 
R17 A2 A2:4 22.2387 
R18 A2:5 A2:4 23.7128 
R19 A2:4 M28:GATE 111.3 
CC47945 A2:4 M11:SRC 2.179e-17
CC48133 A2:4 M28:SRC 4.11e-18
CC48139 M28:GATE N_9:3 6.84e-18
CC48125 M28:GATE M28:SRC 2.514e-17
R20 M11:GATE A2:5 81.5607 
R21 A2 A2:5 22.4407 
R22 A2:6 A2:5 26.843 
R23 A2:5 M27:GATE 111.3 
CC47926 A2:5 ZN:3 1.58e-18
CC47946 A2:5 M11:SRC 2.892e-17
CC48175 A2:5 M26:SRC 4.03e-18
CC48168 M27:GATE M26:SRC 2.572e-17
CC48140 M27:GATE N_9:3 5.96e-18
R24 M9:GATE M25:GATE 738.467 
R25 M25:GATE A2:6 154.179 
CC48183 M25:GATE M24:SRC 4.78e-17
CC48059 M25:GATE N_9:2 2.04e-18
CC48045 M25:GATE N_9:1 3.66e-18
CC48142 M25:GATE N_9:3 4.14e-18
R26 M10:GATE A2:6 94.0755 
R27 M9:GATE A2:6 130.318 
R28 A2:6 M26:GATE 111.3 
CC47932 A2:6 M15:SRC 1.428e-17
CC47937 A2:6 M13:SRC 1.412e-17
CC47922 A2:6 ZN:3 1.978e-17
CC47949 A2:6 M9:SRC 7.412e-17
CC47943 A2:6 M11:SRC 1.48e-17
CC48159 A2:6 N_9:3 1.802e-17
CC48174 A2:6 M26:SRC 1.778e-17
CC48119 A2:6 M30:SRC 1.426e-17
CC48130 A2:6 M28:SRC 1.427e-17
CC48169 M26:GATE M26:SRC 2.67e-17
CC48058 M26:GATE N_9:2 1.61e-18
CC48141 M26:GATE N_9:3 7.37e-18
CC47935 A2 M13:SRC 3.78e-18
CC47920 A2 ZN:3 9.724e-17
CC47942 A2 M11:SRC 3.65e-18
CC48156 A2 N_9:3 7.104e-17
CC48173 A2 M26:SRC 1.14e-18
CC48117 A2 M30:SRC 1.63e-18
CC48129 A2 M28:SRC 1.36e-18
CC47934 M14:GATE M13:SRC 8.48e-18
CC47914 M14:GATE ZN:3 3.49e-18
CC47919 M9:GATE ZN:3 3.3e-18
CC47918 M10:GATE ZN:3 2.8e-18
CC47917 M11:GATE ZN:3 2.84e-18
CC47916 M12:GATE ZN:3 3.74e-18
CC47941 M12:GATE M11:SRC 7.43e-18
CC47913 M15:GATE ZN:3 3.42e-18
CC48113 M30:GATE M30:SRC 2.45e-17
CC48137 M30:GATE N_9:3 6.84e-18
CC48177 M32:GATE M32:SRC 5.103e-17
CC48135 M32:GATE N_9:3 6.4e-18
CC48138 M29:GATE N_9:3 5.89e-18
CC48124 M29:GATE M28:SRC 2.573e-17
C29 A2:3 0 1.402e-17
C30 A2:2 0 2.249e-17
C31 M31:GATE 0 6.316e-17
C32 A2:1 0 5.472e-17
C33 M16:GATE 0 3.09e-17
C34 A2:4 0 2.207e-17
C35 M28:GATE 0 6.277e-17
C36 A2:5 0 1.59e-18
C37 M27:GATE 0 6.453e-17
C38 M25:GATE 0 6.141e-17
C39 A2:6 0 8.665e-17
C40 M26:GATE 0 5.562e-17
C41 A2 0 2.359e-17
C42 M14:GATE 0 4.27e-17
C43 M9:GATE 0 6.479e-17
C44 M10:GATE 0 4.824e-17
C45 M11:GATE 0 3.513e-17
C46 M12:GATE 0 3.246e-17
C47 M13:GATE 0 5.07e-17
C48 M15:GATE 0 5.284e-17
C49 M30:GATE 0 7.374e-17
C50 M32:GATE 0 5.104e-17
C51 M29:GATE 0 6.211e-17
R52 M18:DRN M17:SRC 0.001 
R53 ZN M17:SRC 45.3709 
R54 M17:SRC ZN:1 94.9136 
CC48070 M17:SRC N_9:2 5.47e-18
CC47953 M17:SRC A1:1 1.09e-18
CC48001 M17:SRC A1:4 1.311e-17
CC47995 M17:SRC M17:GATE 2.77e-17
CC47992 M17:SRC M18:GATE 2.689e-17
R55 M21:SRC ZN:1 29.9999 
R56 M19:SRC ZN:1 94.1018 
R57 M23:SRC ZN:1 30.4612 
R58 ZN:1 ZN 0.48933 
CC48016 ZN:1 A1 3.7e-17
CC48007 ZN:1 A1:4 2.43e-17
CC48028 ZN:1 M3:GATE 1.2e-18
CC48039 ZN:1 M23:GATE 8.45e-18
CC48035 ZN:1 M24:GATE 2.95e-18
CC48050 ZN:1 N_9:1 1.3497e-16
CC48075 ZN:1 N_9:2 2.757e-17
CC48085 ZN:1 M22:SRC 7.19e-18
CC48094 ZN:1 M20:SRC 7.43e-18
CC48102 ZN:1 M18:SRC 7.43e-18
CC48108 ZN:1 M17:DRN 1.09e-18
CC47980 ZN:1 M21:GATE 8.49e-18
CC47967 ZN:1 M22:GATE 8.04e-18
CC47996 ZN:1 M17:GATE 3.02e-18
CC47994 ZN:1 M18:GATE 1.126e-17
CC47985 ZN:1 M20:GATE 8.8e-18
CC47989 ZN:1 M19:GATE 7.89e-18
CC47956 ZN:1 A1:1 1.11e-18
CC47963 ZN:1 A1:2 4.2e-18
CC48165 ZN:1 N_9:3 1.646e-17
R59 M19:SRC ZN 44.4938 
R60 ZN ZN:3 0.12133 
CC48015 ZN A1 1.512e-17
CC48006 ZN A1:4 1.94e-17
CC48072 ZN N_9:2 1.05e-18
CC48092 ZN M20:SRC 1.78e-18
CC47984 ZN M20:GATE 3.33e-18
CC47979 ZN M21:GATE 1.68e-18
CC47988 ZN M19:GATE 1.89e-18
R61 M7:SRC ZN:3 71.88 
R62 ZN:2 ZN:3 1.7509 
R63 M3:SRC ZN:3 29.9999 
R64 M5:SRC ZN:3 35.5078 
R65 ZN:3 M1:SRC 30.4724 
CC48008 ZN:3 A1:4 1.638e-17
CC48017 ZN:3 A1 8.087e-17
CC48041 ZN:3 M8:GATE 3.98e-18
CC48042 ZN:3 M7:GATE 2.98e-18
CC48033 ZN:3 M1:GATE 1.98e-18
CC48051 ZN:3 N_9:1 1.79e-18
CC48030 ZN:3 M2:GATE 3.26e-18
CC48029 ZN:3 M3:GATE 5.18e-18
CC48022 ZN:3 M5:GATE 2.87e-18
CC48019 ZN:3 M6:GATE 3.6e-18
CC48025 ZN:3 M4:GATE 3.26e-18
CC47990 ZN:3 M19:GATE 2.58e-18
CC47964 ZN:3 A1:2 1.83e-18
CC47957 ZN:3 A1:1 3.69e-18
CC48166 ZN:3 N_9:3 2.406e-17
R66 M1:SRC M2:DRN 0.001 
CC48005 M1:SRC A1:4 1.539e-17
CC48032 M1:SRC M2:GATE 2.098e-17
CC47955 M1:SRC A1:1 3.758e-17
R67 ZN:2 M5:SRC 207.654 
R68 M5:SRC M6:DRN 0.001 
CC48013 M5:SRC A1 2.66e-18
CC48003 M5:SRC A1:4 1.431e-17
CC48020 M5:SRC M5:GATE 3.98e-18
CC48018 M5:SRC M6:GATE 5.2e-18
CC47972 M5:SRC A1:3 3.36e-17
CC47960 M5:SRC A1:2 1.576e-17
R69 M23:SRC M24:DRN 0.001 
CC48009 M23:SRC A1 1.55e-18
CC48036 M23:SRC M23:GATE 2.783e-17
CC48034 M23:SRC M24:GATE 2.773e-17
CC48047 M23:SRC N_9:1 4.99e-18
CC48061 M23:SRC N_9:2 4.51e-18
CC47998 M23:SRC A1:4 1.3e-17
R70 M3:SRC M4:DRN 0.001 
CC48004 M3:SRC A1:4 1.562e-17
CC48023 M3:SRC M4:GATE 2.088e-17
CC47961 M3:SRC A1:2 2.706e-17
CC47954 M3:SRC A1:1 9.33e-18
R71 M16:SRC M15:SRC 0.001 
R72 M13:SRC M15:SRC 711.195 
R73 M11:SRC M15:SRC 1468.16 
R74 M15:SRC ZN:2 34.3868 
R75 M13:SRC ZN:2 33.5693 
R76 M7:SRC ZN:2 52.7361 
R77 M9:SRC ZN:2 29.9999 
R78 ZN:2 M11:SRC 32.0274 
R79 M13:SRC M11:SRC 1433.26 
R80 M11:SRC M12:DRN 0.001 
R81 M19:SRC M20:DRN 0.001 
CC48067 M19:SRC N_9:2 4.81e-18
CC47983 M19:SRC M20:GATE 2.706e-17
CC48000 M19:SRC A1:4 1.301e-17
CC47986 M19:SRC M19:GATE 2.729e-17
R82 M21:SRC M22:DRN 0.001 
CC48010 M21:SRC A1 1.04e-18
CC48064 M21:SRC N_9:2 4.81e-18
CC47976 M21:SRC M21:GATE 2.748e-17
CC47969 M21:SRC A1:3 1.1e-18
CC47966 M21:SRC M22:GATE 2.82e-17
CC47999 M21:SRC A1:4 1.307e-17
R83 M9:SRC M10:DRN 0.001 
R84 M7:SRC M8:DRN 0.001 
CC48012 M7:SRC A1 7.83e-18
CC48040 M7:SRC M8:GATE 2.439e-17
CC48002 M7:SRC A1:4 4.255e-17
R85 M13:SRC M14:DRN 0.001 
C86 M17:SRC 0 1.232e-17
C87 ZN:1 0 8.3e-18
C88 ZN:3 0 4.2611e-16
C89 M1:SRC 0 4.87e-18
C90 M5:SRC 0 5.38e-18
C91 M23:SRC 0 1.12e-18
C92 M3:SRC 0 6.72e-18
C93 M15:SRC 0 6.69e-18
C94 ZN:2 0 1.652e-17
C95 M11:SRC 0 5.4e-18
C96 M19:SRC 0 2.59e-18
C97 M21:SRC 0 1.81e-18
C98 M9:SRC 0 4.13e-18
C99 M7:SRC 0 7.92e-18
C100 M13:SRC 0 1.006e-17
R101 M3:GATE M19:GATE 1066.52 
R102 A1:1 M19:GATE 275.689 
R103 M19:GATE A1:2 275.689 
CC48097 M19:GATE M18:SRC 2.909e-17
CC48068 M19:GATE N_9:2 7.29e-18
R104 M5:GATE A1:2 247.656 
R105 M4:GATE A1:2 94.0755 
R106 M3:GATE A1:2 233.022 
R107 M20:GATE A1:2 111.3 
R108 A1:1 A1:2 60.2341 
R109 A1:3 A1:2 55.3995 
R110 A1:2 M21:GATE 293 
R111 M5:GATE M21:GATE 1133.5 
R112 M21:GATE A1:3 253.558 
CC48088 M21:GATE M20:SRC 2.938e-17
CC48065 M21:GATE N_9:2 6.39e-18
R113 M6:GATE A1:3 81.9458 
R114 M5:GATE A1:3 214.316 
R115 M22:GATE A1:3 111.3 
R116 A1:4 A1:3 23.7076 
R117 A1:3 A1 22.4649 
R118 M24:GATE A1 237.259 
R119 M8:GATE A1 195.465 
R120 A1 A1:4 16.0695 
CC48048 A1 N_9:1 3.19e-18
CC48157 A1 N_9:3 1.173e-17
CC48189 A1 M24:SRC 1.22e-18
R121 M7:GATE A1:4 81.2035 
R122 M23:GATE A1:4 88.7752 
R123 M24:GATE A1:4 256.16 
R124 A1:4 M8:GATE 211.037 
CC48049 A1:4 N_9:1 2.03e-18
CC48093 A1:4 M20:SRC 5.3e-18
CC48084 A1:4 M22:SRC 5.33e-18
CC48101 A1:4 M18:SRC 5.39e-18
R125 M8:GATE M24:GATE 865.248 
CC48060 M24:GATE N_9:2 5.76e-18
CC48143 M24:GATE N_9:3 1.43e-18
CC48184 M24:GATE M24:SRC 4.737e-17
R126 M1:GATE M17:GATE 635.948 
R127 M17:GATE A1:1 164.389 
CC48105 M17:GATE M17:DRN 5.07e-17
CC48071 M17:GATE N_9:2 9.99e-18
R128 M2:GATE A1:1 94.0755 
R129 M3:GATE A1:1 233.022 
R130 M1:GATE A1:1 138.947 
R131 A1:1 M18:GATE 111.3 
CC48098 M18:GATE M18:SRC 2.938e-17
CC48069 M18:GATE N_9:2 7.26e-18
CC48080 M22:GATE M22:SRC 2.965e-17
CC48063 M22:GATE N_9:2 6.73e-18
CC48089 M20:GATE M20:SRC 2.938e-17
CC48066 M20:GATE N_9:2 6.73e-18
CC48062 M23:GATE N_9:2 6.29e-18
CC48079 M23:GATE M22:SRC 2.954e-17
C132 M19:GATE 0 2.455e-17
C133 A1:2 0 3.498e-17
C134 M21:GATE 0 2.661e-17
C135 A1:3 0 2.989e-17
C136 A1 0 4.695e-17
C137 A1:4 0 7.642e-17
C138 M8:GATE 0 3.317e-17
C139 M24:GATE 0 3.881e-17
C140 M17:GATE 0 2.511e-17
C141 A1:1 0 5.568e-17
C142 M18:GATE 0 1.632e-17
C143 M22:GATE 0 2.629e-17
C144 M20:GATE 0 1.842e-17
C145 M23:GATE 0 3.892e-17
C146 M1:GATE 0 6.427e-17
C147 M7:GATE 0 5.494e-17
C148 M3:GATE 0 5.689e-17
C149 M4:GATE 0 3.187e-17
C150 M5:GATE 0 4.412e-17
C151 M2:GATE 0 2.651e-17
C152 M6:GATE 0 3.994e-17
R153 M26:SRC N_9:1 29.9999 
R154 M28:SRC N_9:1 46.5409 
R155 M22:SRC N_9:1 114.412 
R156 N_9:2 N_9:1 2.37892 
R157 M24:SRC N_9:1 23.6049 
R158 N_9:3 N_9:1 1.70821 
R159 N_9:1 M30:SRC 99.48 
R160 M30:SRC N_9:3 43.6844 
R161 M28:SRC N_9:3 88.9583 
R162 N_9:3 M32:SRC 15.0745 
R163 M24:SRC N_9:2 44.3544 
R164 M17:DRN N_9:2 16.6558 
R165 M18:SRC N_9:2 31.8151 
R166 M20:SRC N_9:2 29.9999 
R167 N_9:2 M22:SRC 42.3141 
R168 M18:SRC M17:DRN 801.044 
C169 N_9:1 0 7.437e-17
C170 M30:SRC 0 4.41e-18
C171 N_9:3 0 1.9275e-16
C172 M32:SRC 0 2.3e-17
C173 M24:SRC 0 1.57e-17
C174 N_9:2 0 1.2682e-16
C175 M22:SRC 0 9.16e-18
C176 M28:SRC 0 4.07e-18
C177 M26:SRC 0 1.37e-17
C178 M20:SRC 0 5.37e-18
C179 M18:SRC 0 1.568e-17
C180 M17:DRN 0 1.815e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
