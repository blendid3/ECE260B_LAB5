.SUBCKT AOI21D2 A1 A2 B ZN
MMM10 M10:DRN M10:GATE M10:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.6e-07  SB=9.4e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 M10:SRC M11:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=4e-07  SB=1.2e-06  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.567  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=8.3e-14  AS=4.7e-14  PD=1.36e-06  PS=7e-07  SA=1.6e-07  SB=1.44e-06  NRD=0.532  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M1:SRC M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.18e-06  SB=4.2e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.2e-07  SB=6.8e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M3:SRC M4:GATE M4:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.6e-07  SB=9.4e-07  NRD=4.12  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=4e-07  SB=1.2e-06  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 vss M6:GATE M6:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=6.2e-14  PD=5.7e-07  PS=1.1e-06  SA=1.6e-07  SB=1.44e-06  NRD=7.648  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 M7:DRN M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.532  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE M8:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.18e-06  SB=4.2e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 M8:SRC M9:GATE M9:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.2e-07  SB=6.8e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
CC90820 M1:SRC A1 1.02e-18
CC90819 M3:SRC A1 1.02e-18
R0 M7:SRC ZN 33.1457 
R1 M6:SRC ZN 30.9965 
R2 M9:SRC ZN 32.2128 
R3 M4:SRC ZN 31.0514 
R4 ZN M1:DRN 32.3409 
CC90826 ZN B:1 1.577e-17
CC90832 ZN M12:GATE 2.74e-18
CC90838 ZN M11:GATE 1.654e-17
CC90801 ZN M12:DRN 1.5e-18
CC90802 ZN M10:SRC 2.354e-17
CC90803 ZN M10:GATE 6.21e-18
CC90804 ZN M8:SRC 3.865e-17
CC90805 ZN M7:GATE 1.35e-18
CC90806 ZN M7:DRN 9.444e-17
CC90807 ZN M4:GATE 8.9e-18
CC90808 ZN M1:GATE 4.86e-18
CC90809 ZN A1 1.5719e-16
CC90842 ZN B 6.911e-17
CC90846 ZN M5:GATE 4.27e-18
CC90856 ZN A2:1 6.33e-18
CC90864 ZN M9:GATE 4.96e-18
CC90873 ZN M8:GATE 5.31e-18
CC90879 ZN A2 4.018e-17
CC90881 ZN M2:GATE 3.08e-18
R5 M1:DRN M4:SRC 1627.46 
CC90818 M1:DRN A1 3.166e-17
R6 M4:SRC M5:DRN 0.001 
CC90825 M4:SRC B:1 2.486e-17
CC90814 M4:SRC A1 3.118e-17
CC90844 M4:SRC M5:GATE 5.08e-18
R7 M7:SRC M9:SRC 886.123 
R8 M9:SRC M10:DRN 0.001 
CC90799 M9:SRC M8:SRC 6.68e-18
CC90800 M9:SRC A1 7.6e-18
CC90860 M9:SRC M9:GATE 2.761e-17
CC90798 M9:SRC M10:GATE 2.942e-17
CC90824 M6:SRC B:1 3.028e-17
CC90841 M6:SRC B 2.95e-18
R9 M7:SRC M8:DRN 0.001 
CC90870 M7:SRC M8:GATE 2.75e-17
CC90792 M7:SRC M8:SRC 6.53e-18
CC90793 M7:SRC M7:GATE 2.775e-17
CC90795 M7:SRC M1:GATE 1.66e-18
CC90796 M7:SRC A1 8.3e-18
C10 ZN 0 1.1235e-16
C11 M1:DRN 0 1.351e-17
C12 M4:SRC 0 6.84e-18
C13 M9:SRC 0 5.97e-18
C14 M6:SRC 0 2.223e-17
C15 M7:SRC 0 5.98e-18
R16 M1:GATE M7:GATE 519.013 
R17 M7:GATE A1 150.526 
CC90853 M7:GATE A2:1 1.083e-17
CC90871 M7:GATE M8:GATE 7.04e-18
CC90787 M7:GATE M7:DRN 2.774e-17
CC90786 M7:GATE M8:SRC 4.32e-18
CC90785 M7:GATE M12:DRN 4.51e-18
R18 M1:GATE A1 124.184 
R19 M4:GATE A1 121.354 
R20 A1 M10:GATE 147.094 
CC90857 A1 A2:1 9.76e-18
CC90843 A1 B 2.18e-18
CC90839 A1 M11:GATE 1.06e-18
CC90827 A1 B:1 7.7e-18
CC90865 A1 M9:GATE 6.28e-18
CC90874 A1 M8:GATE 8.33e-18
CC90880 A1 A2 7.07e-17
CC90885 A1 M3:GATE 3.4e-18
CC90790 A1 M8:SRC 4.39e-18
CC90788 A1 M12:DRN 1.174e-17
CC90791 A1 M7:DRN 1.42e-18
R21 M10:GATE M4:GATE 542.94 
CC90859 M10:GATE M9:GATE 6.89e-18
CC90849 M10:GATE A2:1 4.63e-18
CC90823 M10:GATE B:1 5.93e-18
CC90835 M10:GATE M11:GATE 6.46e-18
CC90783 M10:GATE M10:SRC 2.923e-17
CC90784 M10:GATE M8:SRC 6.84e-18
CC90855 M4:GATE A2:1 1.363e-17
CC90845 M4:GATE M5:GATE 4.03e-18
CC90886 M4:GATE M3:GATE 4.03e-18
CC90878 M1:GATE A2 9.42e-18
CC90883 M1:GATE M2:GATE 1.031e-17
C22 M7:GATE 0 3.693e-17
C23 A1 0 2.293e-17
C24 M10:GATE 0 3.689e-17
C25 M4:GATE 0 3.235e-17
C26 M1:GATE 0 3.495e-17
R27 M12:DRN M8:SRC 124.277 
R28 M7:DRN M8:SRC 118.721 
R29 M8:SRC M10:SRC 121.429 
CC90861 M8:SRC M9:GATE 3.584e-17
CC90851 M8:SRC A2:1 1.13e-17
CC90869 M8:SRC M8:GATE 3.447e-17
CC90837 M8:SRC M11:GATE 7.64e-18
CC90831 M8:SRC M12:GATE 8.39e-18
R30 M12:DRN M10:SRC 118.617 
R31 M10:SRC M7:DRN 124.39 
CC90834 M10:SRC M11:GATE 2.927e-17
R32 M7:DRN M12:DRN 127.308 
CC90866 M12:DRN M8:GATE 1.66e-18
CC90840 M12:DRN B 1.628e-17
CC90828 M12:DRN M12:GATE 2.798e-17
C33 M8:SRC 0 6.48e-18
C34 M10:SRC 0 8.765e-17
C35 M7:DRN 0 2.822e-17
C36 M12:DRN 0 8.783e-17
R37 M12:GATE B:1 111.3 
R38 M6:GATE B:1 83.3024 
R39 B B:1 22 
R40 M5:GATE B:1 130.664 
R41 B:1 M11:GATE 154.587 
R42 M11:GATE M5:GATE 733.433 
C43 M12:GATE 0 4.901e-17
C44 B:1 0 2.943e-17
C45 M11:GATE 0 4.741e-17
C46 M5:GATE 0 4.177e-17
C47 B 0 1.399e-17
C48 M6:GATE 0 4.578e-17
R49 M9:GATE A2:1 111.3 
R50 M3:GATE A2:1 94.0755 
R51 M2:GATE A2:1 201.322 
R52 A2 A2:1 37.7348 
R53 A2:1 M8:GATE 238.184 
R54 M2:GATE M8:GATE 722.167 
R55 M8:GATE A2 448.204 
R56 A2 M2:GATE 378.839 
C57 M9:GATE 0 4.056e-17
C58 A2:1 0 5.278e-17
C59 M8:GATE 0 3.842e-17
C60 A2 0 8.17e-18
C61 M2:GATE 0 5.114e-17
C62 M3:GATE 0 5.648e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
