.SUBCKT LHQD2 D E Q
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=2.68e-07  AD=4.4e-14  AS=3.2e-14  PD=8.6e-07  PS=5.85e-07  SA=1.7e-07  SB=2.34e-07  NRD=0.737  NRS=0.726  SCA=5.723  SCB=0.006  SCC=0.0001074 
MMM11 M11:DRN M11:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=5e-14  AS=3.2e-14  PD=9.4e-07  PS=5.85e-07  SA=2.33e-07  SB=1.88e-07  NRD=0.811  NRS=0.726  SCA=11.263  SCB=0.013  SCC=0.0008706 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=2.67e-07  AD=4e-14  AS=1.8e-14  PD=8.3e-07  PS=4e-07  SA=1.55e-07  SB=6.18e-07  NRD=1.392  NRS=19.974  SCA=6.917  SCB=0.007  SCC=0.000196 
MMM12 vdd M12:GATE M12:SRC vdd pch L=6e-08 W=3.44e-07  AD=5.3e-14  AS=2.4e-14  PD=9.9e-07  PS=4.8e-07  SA=1.55e-07  SB=4.87e-07  NRD=1.424  NRS=21.508  SCA=12.895  SCB=0.014  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=1.58e-07  AD=1.5e-14  AS=1e-14  PD=3.5e-07  PS=2.9e-07  SA=8.45e-07  SB=4.35e-07  NRD=10.929  NRS=34.621  SCA=6.231  SCB=0.006  SCC=0.0001038 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=1.5e-07  AD=1.5e-14  AS=1e-14  PD=3.5e-07  PS=2.9e-07  SA=8.45e-07  SB=4.35e-07  NRD=6.977  NRS=48.752  SCA=6.744  SCB=0.007  SCC=0.0001603 
MMM3 M1:SRC M3:GATE M3:SRC vss nch L=6.1e-08 W=2.6e-07  AD=1.8e-14  AS=3.4e-14  PD=4e-07  PS=6.21e-07  SA=3.55e-07  SB=3.45e-07  NRD=19.974  NRS=4.774  SCA=6.917  SCB=0.007  SCC=0.000196 
MMM14 M14:DRN M14:GATE vdd vdd pch L=6e-08 W=1.5e-07  AD=2.6e-14  AS=1.5e-14  PD=6.5e-07  PS=3.5e-07  SA=1.115e-06  SB=1.75e-07  NRD=1.195  NRS=6.977  SCA=6.744  SCB=0.007  SCC=0.0001603 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=1.58e-07  AD=2.6e-14  AS=1.5e-14  PD=6.5e-07  PS=3.5e-07  SA=1.115e-06  SB=1.75e-07  NRD=1.195  NRS=10.929  SCA=6.231  SCB=0.006  SCC=0.0001038 
MMM15 M13:SRC M15:GATE M15:SRC vdd pch L=6e-08 W=1.51e-07  AD=1e-14  AS=1.8e-14  PD=2.9e-07  PS=3.49e-07  SA=6.45e-07  SB=6.35e-07  NRD=48.752  NRS=0.812  SCA=6.744  SCB=0.007  SCC=0.0001603 
MMM5 M2:SRC M5:GATE M3:SRC vss nch L=6e-08 W=1.58e-07  AD=1e-14  AS=2e-14  PD=2.9e-07  PS=3.59e-07  SA=6.45e-07  SB=6.35e-07  NRD=34.621  NRS=0.881  SCA=6.231  SCB=0.006  SCC=0.0001038 
MMM16 M15:SRC M16:GATE M12:SRC vdd pch L=6e-08 W=3.4e-07  AD=4.1e-14  AS=2.4e-14  PD=7.91e-07  PS=4.8e-07  SA=3.55e-07  SB=2.23e-07  NRD=11.184  NRS=21.508  SCA=12.895  SCB=0.014  SCC=0.001 
MMM6 vss M6:GATE M6:SRC vss nch L=6e-08 W=3.97e-07  AD=5.1e-14  AS=3.9e-14  PD=1.04e-06  PS=5.9e-07  SA=3.9e-07  SB=1.3e-07  NRD=1.615  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 vdd M17:GATE M17:SRC vdd pch L=6e-08 W=5.24e-07  AD=6.8e-14  AS=5.2e-14  PD=1.3e-06  PS=7.2e-07  SA=3.91e-07  SB=1.3e-07  NRD=1.865  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 M7:DRN M7:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=5.1e-14  PD=5.9e-07  PS=1.04e-06  SA=1.3e-07  SB=3.9e-07  NRD=4.183  NRS=1.615  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M18:DRN M18:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.8e-14  PD=7.2e-07  PS=1.3e-06  SA=1.3e-07  SB=3.9e-07  NRD=2.057  NRS=1.865  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=2.02e-07  AD=3.4e-14  AS=2e-14  PD=7.4e-07  PS=3.95e-07  SA=1.75e-07  SB=4.7e-07  NRD=0.947  NRS=8.494  SCA=18.109  SCB=0.02  SCC=0.002 
MMM9 M9:DRN M9:GATE vss vss nch L=6e-08 W=2.02e-07  AD=4.1e-14  AS=2e-14  PD=8.1e-07  PS=3.95e-07  SA=4.35e-07  SB=2.1e-07  NRD=1.119  NRS=8.494  SCA=18.109  SCB=0.02  SCC=0.002 
R0 Q M7:DRN 15.2336 
R1 M7:DRN M6:SRC 0.001 
CC86309 M7:DRN M7:GATE 8.19e-18
CC86266 M7:DRN N_26:1 1.481e-17
CC86273 M7:DRN N_26:2 7.659e-17
CC86221 M7:DRN M4:DRN 1.92e-18
CC86314 M7:DRN M6:GATE 1.628e-17
R2 Q M18:DRN 15.3641 
CC86285 Q M18:GATE 7.59e-18
CC86308 Q M4:GATE 1.722e-17
CC86289 Q M17:GATE 2.695e-17
CC86217 Q M14:DRN 5.951e-17
CC86271 Q N_26:1 1.05e-18
CC86276 Q N_26:2 4.26e-18
CC86316 Q M6:GATE 1.468e-17
CC86313 Q M7:GATE 3.89e-18
R3 M18:DRN M17:SRC 0.001 
CC86220 M18:DRN M4:DRN 1.43e-18
CC86286 M18:DRN M17:GATE 4.735e-17
CC86290 M18:DRN M14:GATE 6.44e-18
CC86258 M18:DRN N_26:1 7.22e-18
CC86277 M18:DRN M18:GATE 4.776e-17
C4 M7:DRN 0 2.67e-18
C5 Q 0 9.053e-17
C6 M18:DRN 0 6.9e-18
R7 E M8:GATE 84.0774 
R8 M8:GATE M10:GATE 396.24 
CC86246 M8:GATE M9:GATE 3.87e-18
CC86253 M8:GATE M8:DRN 3.812e-17
R9 M10:GATE E 170.222 
CC86251 M10:GATE M8:DRN 1.413e-17
CC86231 M10:GATE M11:GATE 9.06e-18
CC86235 M10:GATE M10:DRN 2.962e-17
CC86248 E M9:GATE 5.99e-18
CC86255 E M8:DRN 3.752e-17
CC86233 E M11:GATE 3e-18
CC86237 E M10:DRN 7.681e-17
C10 M8:GATE 0 3.014e-17
C11 M10:GATE 0 5.383e-17
C12 E 0 1.959e-17
R13 M1:GATE D 138.814 
R14 D M12:GATE 114.318 
CC86234 D M11:GATE 2.84e-18
CC86211 D M11:DRN 4.72e-18
CC86212 D M9:DRN 9.24e-18
CC86213 D M3:GATE 1.0095e-16
CC86228 D M16:GATE 7.34e-18
CC86256 D M8:DRN 5.55e-18
R15 M12:GATE M1:GATE 468.183 
CC86209 M12:GATE M11:DRN 2.94e-18
CC86210 M12:GATE M9:DRN 1.389e-17
CC86224 M12:GATE M16:GATE 2.443e-17
CC86214 M1:GATE M11:DRN 2.066e-17
CC86215 M1:GATE M9:DRN 2.19e-18
CC86216 M1:GATE M3:GATE 1.109e-17
C16 D 0 3.074e-17
C17 M12:GATE 0 4.948e-17
C18 M1:GATE 0 2.842e-17
R19 M2:GATE M4:DRN 305.363 
R20 M14:DRN M4:DRN 74.2872 
R21 M4:DRN M13:GATE 384.203 
CC86306 M4:DRN M4:GATE 2.387e-17
CC86296 M4:DRN M14:GATE 3.86e-18
CC86207 M4:DRN M9:DRN 2.55e-18
CC86268 M4:DRN N_26:1 3.547e-17
CC86241 M4:DRN M5:GATE 2.755e-17
CC86310 M4:DRN M7:GATE 9.66e-18
CC86284 M4:DRN M18:GATE 4.92e-18
CC86320 M4:DRN M3:SRC 5.7e-18
CC86274 M4:DRN N_26:2 1.602e-17
R22 M2:GATE M13:GATE 448.316 
R23 M13:GATE M14:DRN 399.419 
CC86300 M13:GATE M15:SRC 2.33e-18
CC86294 M13:GATE M14:GATE 2.31e-18
CC86262 M13:GATE N_26:1 4.935e-17
CC86239 M13:GATE M5:GATE 2.91e-18
CC86204 M13:GATE M9:DRN 9.39e-18
CC86203 M13:GATE M15:GATE 1.151e-17
R24 M14:DRN M2:GATE 317.457 
CC86293 M14:DRN M14:GATE 3.15e-17
CC86261 M14:DRN N_26:1 1.2119e-16
CC86280 M14:DRN M18:GATE 3.72e-18
CC86243 M2:GATE M5:GATE 7.27e-18
CC86307 M2:GATE M4:GATE 6.94e-18
CC86275 M2:GATE N_26:2 1.682e-17
CC86270 M2:GATE N_26:1 3.68e-18
C25 M4:DRN 0 9.685e-17
C26 M13:GATE 0 5.567e-17
C27 M14:DRN 0 1.836e-17
C28 M2:GATE 0 5.895e-17
R29 M15:GATE M9:DRN 227.915 
R30 M11:DRN M9:DRN 83.5527 
R31 M9:DRN M3:GATE 213.019 
CC86245 M9:DRN M9:GATE 5.29e-17
CC86240 M9:DRN M5:GATE 1.258e-17
CC86265 M9:DRN N_26:1 9.18e-18
CC86318 M9:DRN M3:SRC 2.911e-17
CC86252 M9:DRN M8:DRN 2.346e-17
CC86236 M9:DRN M10:DRN 1.629e-17
CC86232 M9:DRN M11:GATE 2.211e-17
CC86301 M9:DRN M15:SRC 2.604e-17
CC86226 M9:DRN M16:GATE 2.234e-17
R32 M15:GATE M3:GATE 527.025 
R33 M3:GATE M11:DRN 218.615 
CC86242 M3:GATE M5:GATE 1.81e-18
CC86269 M3:GATE N_26:1 1.501e-17
CC86321 M3:GATE M3:SRC 3.33e-18
CC86227 M3:GATE M16:GATE 9.19e-18
R34 M11:DRN M15:GATE 233.902 
CC86264 M11:DRN N_26:1 3.961e-17
CC86250 M11:DRN M8:DRN 4.31e-18
CC86230 M11:DRN M11:GATE 1.913e-17
CC86225 M11:DRN M16:GATE 3.17e-18
CC86238 M15:GATE M5:GATE 3.42e-18
CC86260 M15:GATE N_26:1 6.931e-17
CC86299 M15:GATE M15:SRC 1.961e-17
CC86222 M15:GATE M16:GATE 8.79e-18
C35 M9:DRN 0 4.507e-17
C36 M3:GATE 0 1.476e-17
C37 M11:DRN 0 1.9817e-16
C38 M15:GATE 0 3.904e-17
R39 M9:GATE M10:DRN 241.45 
R40 M8:DRN M10:DRN 79.2081 
R41 M10:DRN M11:GATE 326.017 
R42 M9:GATE M11:GATE 239.974 
R43 M8:DRN M11:GATE 323.831 
R44 M11:GATE M16:GATE 433.274 
R45 M16:GATE M5:GATE 270.3 
CC86317 M16:GATE M3:SRC 1.16e-17
CC86298 M16:GATE M15:SRC 2.292e-17
CC86259 M16:GATE N_26:1 1.035e-17
CC86302 M5:GATE M15:SRC 3.51e-18
CC86319 M5:GATE M3:SRC 2.281e-17
CC86267 M5:GATE N_26:1 1.371e-17
R46 M8:DRN M9:GATE 239.833 
C47 M10:DRN 0 5.489e-17
C48 M11:GATE 0 7.921e-17
C49 M16:GATE 0 1.1874e-16
C50 M5:GATE 0 1.327e-17
C51 M8:DRN 0 6.478e-17
C52 M9:GATE 0 1.934e-17
R53 M17:GATE M6:GATE 636.814 
R54 M6:GATE N_26:2 140.812 
R55 M7:GATE N_26:2 95.3999 
R56 M18:GATE N_26:2 109.975 
R57 M17:GATE N_26:2 162.326 
R58 M14:GATE N_26:2 373.501 
R59 M4:GATE N_26:2 358.562 
R60 N_26:2 N_26:1 81.0258 
R61 M14:GATE N_26:1 213.557 
R62 M4:GATE N_26:1 205.013 
R63 M3:SRC N_26:1 30.9055 
R64 N_26:1 M15:SRC 30.495 
R65 M4:GATE M14:GATE 945.038 
C66 M6:GATE 0 3.509e-17
C67 N_26:2 0 1.717e-17
C68 N_26:1 0 8.134e-17
C69 M15:SRC 0 9.99e-18
C70 M3:SRC 0 1.029e-17
C71 M4:GATE 0 1.858e-17
C72 M14:GATE 0 6.455e-17
C73 M17:GATE 0 4.757e-17
C74 M18:GATE 0 4.183e-17
C75 M7:GATE 0 2.929e-17
.ENDS
*.SCALE METER 
.GLOBAL VSS VDD
