.SUBCKT ND2D4 A1 A2 ZN
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.72e-06  SB=4.6e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.46e-06  SB=7.2e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7.8e-14  AS=3.9e-14  PD=1.18e-06  PS=5.9e-07  SA=1.98e-06  SB=2e-07  NRD=0.554  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.2e-06  SB=9.8e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M1:SRC M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.72e-06  SB=4.6e-07  NRD=4.12  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.4e-07  SB=1.24e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.46e-06  SB=7.2e-07  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=1.5e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M3:SRC M4:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.2e-06  SB=9.8e-07  NRD=4.12  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vdd M15:GATE M15:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=1.76e-06  NRD=2.099  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.4e-07  SB=1.24e-06  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=2.02e-06  NRD=2.057  NRS=0.427  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M5:SRC M6:GATE M6:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=1.5e-06  NRD=4.12  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 M7:DRN M7:GATE M7:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=1.76e-06  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M7:SRC M8:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.2e-14  PD=5.9e-07  PS=1.1e-06  SA=1.6e-07  SB=2.02e-06  NRD=4.12  NRS=0.462  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.24e-07  AD=1.04e-13  AS=5.2e-14  PD=1.44e-06  PS=7.2e-07  SA=1.98e-06  SB=2e-07  NRD=1.435  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M5:GATE A2:1 78.6162 
R1 A2 A2:1 22 
R2 M4:GATE A2:1 125.092 
R3 M12:GATE A2:1 147.994 
R4 A2:1 M13:GATE 111.3 
CC45097 A2:1 M14:GATE 1.97e-18
CC45089 A2:1 A1:2 9.81e-18
CC45084 A2:1 A1:1 7.47e-18
CC45114 A2:1 A1 1.113e-17
CC45131 A2:1 M3:GATE 1.9e-18
CC45181 A2:1 ZN 1.75e-18
CC45094 M13:GATE M14:GATE 7.5e-18
CC45079 M13:GATE A1:1 1.78e-18
CC45107 M13:GATE A1 5.25e-18
CC45161 M13:GATE M13:SRC 2.851e-17
CC45170 M13:GATE ZN 2.58e-18
R5 M8:GATE A2:2 77.38 
R6 M1:GATE A2:2 9568.71 
R7 M9:GATE A2:2 11698.8 
R8 A2 A2:2 24.702 
R9 A2:2 M16:GATE 94.6047 
CC45092 A2:2 M15:GATE 1.77e-18
CC45083 A2:2 A1:1 1.641e-17
CC45119 A2:2 M6:GATE 4.78e-18
CC45143 A2:2 ZN:1 1.008e-17
CC45090 M16:GATE M15:GATE 2.98e-18
CC45132 M16:GATE ZN:1 4.64e-18
CC45183 M16:GATE M16:DRN 4.757e-17
CC45167 M16:GATE ZN 1.06e-18
R10 M12:GATE M4:GATE 828.301 
CC45085 M12:GATE A1:2 4e-18
CC45108 M12:GATE A1 6.58e-18
CC45099 M12:GATE M11:GATE 7.85e-18
CC45152 M12:GATE M11:SRC 2.782e-17
CC45171 M12:GATE ZN 2.88e-18
CC45086 M4:GATE A1:2 2.35e-18
CC45110 M4:GATE A1 2.21e-18
CC45128 M4:GATE M3:GATE 4.07e-18
R11 M1:GATE A2 124.52 
R12 A2 M9:GATE 152.239 
CC45088 A2 A1:2 2.478e-17
CC45082 A2 A1:1 4.34e-18
CC45123 A2 M7:GATE 8.39e-18
CC45118 A2 M6:GATE 4.48e-18
CC45112 A2 A1 6.251e-17
CC45105 A2 M10:GATE 2.05e-18
CC45149 A2 M9:SRC 1.05e-18
CC45141 A2 ZN:1 8.018e-17
CC45130 A2 M3:GATE 2.61e-18
CC45126 A2 M2:GATE 6.56e-18
CC45199 A2 M2:SRC 4.6e-18
CC45194 A2 M6:SRC 8.23e-18
CC45186 A2 M16:DRN 1.06e-18
CC45178 A2 ZN 1.2267e-16
R13 M9:GATE M1:GATE 464.211 
CC45103 M9:GATE M10:GATE 7.47e-18
CC45148 M9:GATE M9:SRC 2.802e-17
CC45174 M9:GATE ZN 1.671e-17
CC45087 M1:GATE A1:2 1.103e-17
CC45140 M1:GATE ZN:1 3.34e-18
CC45125 M1:GATE M2:GATE 1.097e-17
CC45177 M1:GATE ZN 1.35e-18
CC45116 M5:GATE M6:GATE 4.52e-18
CC45109 M5:GATE A1 7.28e-18
CC45121 M8:GATE M7:GATE 4.11e-18
C14 A2:1 0 7.79e-17
C15 M13:GATE 0 7.674e-17
C16 A2:2 0 7.517e-17
C17 M16:GATE 0 9.413e-17
C18 M12:GATE 0 7.451e-17
C19 M4:GATE 0 4.438e-17
C20 A2 0 3.4949e-16
C21 M9:GATE 0 8.142e-17
C22 M1:GATE 0 3.983e-17
C23 M5:GATE 0 3.592e-17
C24 M8:GATE 0 4.955e-17
R25 M3:GATE A1:2 80.1627 
CC45175 M3:GATE ZN 2.45e-18
R26 A1 A1:2 23.8488 
R27 M10:GATE A1:2 149.317 
R28 M2:GATE A1:2 126.209 
R29 A1:2 M11:GATE 111.3 
CC45182 A1:2 ZN 1.059e-17
CC45195 A1:2 M2:SRC 7.278e-17
CC45153 M11:GATE M11:SRC 2.867e-17
CC45172 M11:GATE ZN 3.22e-18
R30 M2:GATE M10:GATE 806.639 
CC45176 M2:GATE ZN 5.43e-18
CC45147 M10:GATE M9:SRC 2.819e-17
CC45173 M10:GATE ZN 9.93e-18
R31 M6:GATE A1 220.014 
R32 M14:GATE A1 305.98 
R33 A1 A1:1 47.8744 
CC45179 A1 ZN 1.4655e-16
CC45193 A1 M6:SRC 9.33e-18
CC45142 A1 ZN:1 5.044e-17
CC45156 A1 M11:SRC 7.73e-18
CC45164 A1 M13:SRC 7.01e-18
R34 M7:GATE A1:1 94.0755 
R35 M6:GATE A1:1 172.834 
R36 M14:GATE A1:1 240.366 
R37 A1:1 M15:GATE 111.3 
CC45180 A1:1 ZN 1.15e-18
CC45191 A1:1 M6:SRC 6.423e-17
CC45144 A1:1 ZN:1 1.524e-17
CC45184 M15:GATE M16:DRN 4.757e-17
CC45133 M15:GATE ZN:1 7.49e-18
CC45168 M15:GATE ZN 1.54e-18
R38 M14:GATE M6:GATE 1104.64 
CC45134 M14:GATE ZN:1 2.7e-18
CC45160 M14:GATE M13:SRC 2.802e-17
CC45169 M14:GATE ZN 2.99e-18
CC45139 M6:GATE ZN:1 2.37e-18
CC45138 M7:GATE ZN:1 4.41e-18
C39 M3:GATE 0 3.053e-17
C40 A1:2 0 1.409e-17
C41 M11:GATE 0 7.814e-17
C42 M2:GATE 0 3.671e-17
C43 M10:GATE 0 8.283e-17
C44 A1 0 1.469e-17
C45 A1:1 0 1.441e-17
C46 M15:GATE 0 7.444e-17
C47 M14:GATE 0 8.277e-17
C48 M6:GATE 0 3.586e-17
C49 M7:GATE 0 3.103e-17
R50 ZN:1 M13:SRC 44.0058 
R51 M14:DRN M13:SRC 0.001 
R52 M13:SRC ZN 99.5258 
R53 M9:SRC ZN 30.1165 
R54 ZN:1 ZN 2.48876 
R55 M11:SRC ZN 46.2116 
R56 ZN M2:SRC 31.2148 
R57 M2:SRC M3:DRN 0.001 
R58 M12:DRN M11:SRC 0.001 
R59 M11:SRC ZN:1 92.2588 
R60 M16:DRN ZN:1 15.0625 
R61 ZN:1 M6:SRC 30.8752 
R62 M6:SRC M7:DRN 0.001 
R63 M16:DRN M15:SRC 0.001 
R64 M9:SRC M10:DRN 0.001 
C65 M13:SRC 0 8.82e-18
C66 ZN 0 1.7034e-16
C67 M11:SRC 0 9e-18
C68 ZN:1 0 8.555e-17
C69 M16:DRN 0 6.92e-18
C70 M9:SRC 0 3.24e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
