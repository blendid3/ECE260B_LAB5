.SUBCKT INVD0 I ZN
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=1.95e-07  AD=4.8e-14  AS=3.6e-14  PD=8.8e-07  PS=7.6e-07  SA=1.85e-07  SB=2.45e-07  NRD=1.292  NRS=0.996  SCA=9.847  SCB=0.012  SCC=0.0005443 
MMM2 M2:DRN M2:GATE vdd vdd pch L=6e-08 W=2.6e-07  AD=6e-14  AS=4.4e-14  PD=9.8e-07  PS=8.6e-07  SA=1.7e-07  SB=2.3e-07  NRD=0.946  NRS=0.737  SCA=5.375  SCB=0.005  SCC=8.277e-05 
R0 M1:DRN ZN 30.3572 
CC38067 M1:DRN M1:GATE 2.376e-17
CC38064 M1:DRN I 1.248e-17
R1 ZN M2:DRN 30.5759 
CC38062 ZN M2:GATE 6.71e-18
CC38065 ZN I 6.254e-17
CC38066 ZN M1:GATE 9.65e-18
CC38061 M2:DRN M2:GATE 2.995e-17
CC38063 M2:DRN I 2.88e-18
C2 M1:DRN 0 2.146e-17
C3 ZN 0 1.2015e-16
C4 M2:DRN 0 2.967e-17
R5 M2:GATE I 165.276 
R6 I M1:GATE 115.078 
R7 M1:GATE M2:GATE 584.162 
C8 I 0 8.345e-17
C9 M1:GATE 0 4.325e-17
C10 M2:GATE 0 7.705e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
