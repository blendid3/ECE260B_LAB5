.SUBCKT INVD2 I ZN
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.6e-14  AS=3.9e-14  PD=1.12e-06  PS=5.9e-07  SA=4.3e-07  SB=1.7e-07  NRD=0.583  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=6.6e-14  AS=3.9e-14  PD=1.12e-06  PS=5.9e-07  SA=1.7e-07  SB=4.3e-07  NRD=0.583  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vdd M3:GATE M3:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.8e-14  AS=5.2e-14  PD=1.38e-06  PS=7.2e-07  SA=4.3e-07  SB=1.7e-07  NRD=0.538  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 vdd M4:GATE M4:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.8e-14  AS=5.2e-14  PD=1.38e-06  PS=7.2e-07  SA=1.7e-07  SB=4.25e-07  NRD=0.538  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M4:SRC ZN 15.3743 
R1 ZN M2:SRC 15.2507 
CC38174 ZN I:1 2.013e-17
CC38183 ZN M2:GATE 3.7e-18
CC38176 ZN M4:GATE 4.66e-18
CC38178 ZN M3:GATE 9.39e-18
CC38182 ZN I 4.07e-17
R2 M2:SRC M1:SRC 0.001 
CC38181 M2:SRC I 5.03e-18
CC38173 M2:SRC I:1 7.382e-17
CC38186 M2:SRC M1:GATE 2.003e-17
CC38179 M2:SRC M3:GATE 8.59e-18
CC38184 M2:SRC M2:GATE 8.86e-18
R3 M3:SRC M4:SRC 0.001 
CC38172 M4:SRC I:1 9.31e-18
CC38180 M4:SRC I 6.13e-18
CC38175 M4:SRC M4:GATE 4.599e-17
CC38177 M4:SRC M3:GATE 4.748e-17
C4 ZN 0 1.9977e-16
C5 M2:SRC 0 7.34e-18
C6 M4:SRC 0 1.188e-17
R7 M2:GATE I:1 94.0755 
R8 M1:GATE I:1 138.947 
R9 M3:GATE I:1 164.389 
R10 I I:1 34.6266 
R11 I:1 M4:GATE 111.3 
R12 M3:GATE M1:GATE 635.948 
C13 M2:GATE 0 5.433e-17
C14 I:1 0 4.901e-17
C15 M4:GATE 0 8.136e-17
C16 I 0 7.299e-17
C17 M3:GATE 0 7.597e-17
C18 M1:GATE 0 5.982e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
