.SUBCKT NR2D3 A1 A2 ZN
MMM10 M9:SRC M10:GATE M10:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=9.2e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 M11:DRN M11:GATE M11:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=1.18e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.97e-07  AD=5.5e-14  AS=3.9e-14  PD=1.06e-06  PS=5.9e-07  SA=1.44e-06  SB=1.4e-07  NRD=1.549  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M11:SRC M12:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=1.44e-06  NRD=2.099  NRS=0.532  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=1.18e-06  SB=4e-07  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=9.4e-07  SB=6.4e-07  NRD=7.648  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=9e-07  NRD=4.183  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=1.16e-06  NRD=4.537  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.2e-14  PD=5.9e-07  PS=1.1e-06  SA=1.6e-07  SB=1.42e-06  NRD=4.183  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 M7:DRN M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.532  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M7:SRC M8:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.18e-06  SB=4.2e-07  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=9.4e-07  SB=6.6e-07  NRD=6.61  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
CC47726 M7:SRC A1 1.09e-18
CC47681 M11:SRC A2 1.09e-18
R0 ZN:1 ZN 0.08657 
R1 ZN M10:SRC 30.8391 
CC47708 ZN M11:GATE 4.19e-18
CC47714 ZN M10:GATE 8.67e-18
CC47720 ZN M7:GATE 8.25e-18
CC47733 ZN A1 3.28e-18
CC47676 ZN M9:GATE 7.48e-18
CC47679 ZN M8:GATE 7.25e-18
CC47686 ZN A2 7.139e-17
CC47671 ZN A2:1 2.34e-18
R2 M10:SRC M11:DRN 0.001 
CC47696 M10:SRC A1:1 7.84e-18
CC47706 M10:SRC M11:GATE 2.821e-17
CC47711 M10:SRC M10:GATE 2.766e-17
CC47682 M10:SRC A2 6.24e-18
R3 M6:DRN M5:SRC 0.001 
R4 ZN:1 M5:SRC 35.3795 
R5 M3:SRC M5:SRC 598.375 
R6 M5:SRC M1:SRC 894.751 
CC47699 M5:SRC A1:1 2.641e-17
CC47693 M5:SRC M6:GATE 1.12e-17
CC47745 M5:SRC M5:GATE 2.21e-18
CC47683 M5:SRC A2 2.278e-17
R7 ZN:1 M1:SRC 33.4514 
R8 M3:SRC M1:SRC 877.561 
R9 M1:SRC M2:DRN 0.001 
CC47732 M1:SRC A1 3.659e-17
CC47752 M1:SRC M1:GATE 2.31e-18
CC47689 M1:SRC M2:GATE 2.31e-18
CC47670 M1:SRC A2:1 2.394e-17
CC47685 M1:SRC A2 3.18e-18
R10 ZN:1 M3:SRC 34.6997 
R11 M3:SRC M4:DRN 0.001 
CC47700 M3:SRC A1:1 1.407e-17
CC47729 M3:SRC A1 1.964e-17
CC47739 M3:SRC M4:GATE 2.31e-18
CC47669 M3:SRC A2:1 2.647e-17
CC47691 M3:SRC M3:GATE 2.31e-18
R12 ZN:1 M7:DRN 29.9999 
CC47704 ZN:1 A1:1 5.92e-18
CC47716 ZN:1 M10:GATE 3.34e-18
CC47722 ZN:1 M7:GATE 1.674e-17
CC47694 ZN:1 M6:GATE 3.21e-18
CC47736 ZN:1 A1 1.3622e-16
CC47743 ZN:1 M4:GATE 2.27e-18
CC47749 ZN:1 M5:GATE 5.56e-18
CC47754 ZN:1 M1:GATE 1.302e-17
CC47687 ZN:1 A2 3.493e-17
CC47672 ZN:1 A2:1 9.81e-18
CC47680 ZN:1 M8:GATE 2.88e-18
CC47690 ZN:1 M2:GATE 6.54e-18
CC47719 M7:DRN M7:GATE 2.741e-17
C13 ZN 0 8.834e-17
C14 M10:SRC 0 3.94e-18
C15 M5:SRC 0 1.514e-17
C16 M1:SRC 0 1.407e-17
C17 M3:SRC 0 1.389e-17
C18 ZN:1 0 1.1886e-16
C19 M7:DRN 0 1.795e-17
R20 A2:1 M8:GATE 226.529 
R21 M2:GATE M8:GATE 768.451 
R22 M8:GATE A2 461.037 
CC47718 M8:GATE M7:GATE 1.405e-17
R23 M12:GATE A2 149.226 
R24 M6:GATE A2 119.495 
R25 A2:1 A2 39.9913 
R26 A2 M2:GATE 389.689 
CC47753 A2 M1:GATE 4.87e-18
CC47734 A2 A1 1.008e-16
CC47709 A2 M11:GATE 9.7e-18
CC47715 A2 M10:GATE 8.93e-18
CC47702 A2 A1:1 9.75e-18
R27 M2:GATE A2:1 191.47 
CC47751 M2:GATE M1:GATE 3.21e-18
CC47731 M2:GATE A1 5.86e-18
R28 M9:GATE A2:1 111.3 
R29 A2:1 M3:GATE 94.0755 
CC47735 A2:1 A1 2.057e-17
CC47742 A2:1 M4:GATE 3.16e-18
CC47703 A2:1 A1:1 6.27e-18
CC47730 M3:GATE A1 6e-18
CC47740 M3:GATE M4:GATE 3.29e-18
CC47697 M9:GATE A1:1 1.59e-18
CC47712 M9:GATE M10:GATE 1.347e-17
R30 M6:GATE M12:GATE 541.822 
CC47744 M6:GATE M5:GATE 3.09e-18
CC47698 M6:GATE A1:1 2.05e-18
CC47695 M12:GATE A1:1 1.352e-17
CC47705 M12:GATE M11:GATE 1.439e-17
C31 M8:GATE 0 6.064e-17
C32 A2 0 9.321e-17
C33 M2:GATE 0 3.6e-17
C34 A2:1 0 1.848e-17
C35 M3:GATE 0 3.638e-17
C36 M9:GATE 0 5.54e-17
C37 M6:GATE 0 5.037e-17
C38 M12:GATE 0 8.694e-17
R39 M5:GATE A1:1 94.0755 
R40 M4:GATE A1:1 201.305 
R41 M10:GATE A1:1 270.554 
R42 A1 A1:1 53.4785 
R43 A1:1 M11:GATE 111.3 
R44 A1 M7:GATE 150.491 
R45 M7:GATE M1:GATE 519.241 
R46 M1:GATE A1 124.156 
R47 M4:GATE A1 205.874 
R48 A1 M10:GATE 276.694 
R49 M10:GATE M4:GATE 1041.53 
C50 M5:GATE 0 4.386e-17
C51 A1:1 0 1.48e-17
C52 M11:GATE 0 3.7e-17
C53 M7:GATE 0 4.589e-17
C54 M1:GATE 0 3.758e-17
C55 A1 0 1.622e-17
C56 M10:GATE 0 4.487e-17
C57 M4:GATE 0 4.154e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
