.SUBCKT AOI21D4 A1 A2 B ZN
MMM20 M19:SRC M20:GATE M20:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.225e-06  SB=9.37e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 M21:DRN M21:GATE M21:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.65e-07  SB=1.197e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M21:SRC M22:GATE M22:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7.05e-07  SB=1.457e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 M23:DRN M23:GATE M23:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.45e-07  SB=1.735e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 M23:SRC M24:GATE M24:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=9.6e-14  PD=7.2e-07  PS=1.41e-06  SA=1.85e-07  SB=1.995e-06  NRD=2.099  NRS=0.549  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE M10:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.05e-07  SB=4.17e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 M10:SRC M11:GATE M11:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.45e-07  SB=6.7e-07  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.93e-06  SB=1.6e-07  NRD=0.462  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE M12:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=7.2e-14  PD=5.9e-07  PS=1.15e-06  SA=1.85e-07  SB=9.37e-07  NRD=4.183  NRS=0.609  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=1.67e-06  SB=4.2e-07  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=8.9e-07  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=1.43e-06  SB=6.6e-07  NRD=7.648  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M13:SRC M14:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=6.3e-07  SB=4.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4.3e-14  PD=5.9e-07  PS=6.1e-07  SA=1.17e-06  SB=9.2e-07  NRD=4.183  NRS=1.112  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vdd M15:GATE M15:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=3.9e-07  SB=6.6e-07  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.9e-07  AD=4.3e-14  AS=3.9e-14  PD=6.1e-07  PS=5.9e-07  SA=8.9e-07  SB=1.2e-06  NRD=1.112  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M15:SRC M16:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.8e-14  PD=7.2e-07  PS=1.3e-06  SA=1.3e-07  SB=9.2e-07  NRD=2.057  NRS=1.865  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M5:SRC M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=6.3e-07  SB=1.46e-06  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 M17:DRN M17:GATE M17:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.1e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.995e-06  SB=1.57e-07  NRD=0.53  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=3.9e-07  SB=1.7e-06  NRD=7.648  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M17:SRC M18:GATE M18:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.735e-06  SB=4.17e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M7:SRC M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=5.1e-14  PD=5.9e-07  PS=1.04e-06  SA=1.3e-07  SB=1.96e-06  NRD=4.183  NRS=1.615  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 M19:DRN M19:GATE M19:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.475e-06  SB=6.77e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 M9:DRN M9:GATE M9:SRC vss nch L=6e-08 W=3.9e-07  AD=6.1e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=9.65e-07  SB=1.57e-07  NRD=0.562  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
R0 M7:SRC N_11:1 29.9999 
R1 M5:SRC N_11:1 30.5338 
R2 M10:SRC N_11:1 33.0021 
R3 M9:DRN N_11:1 31.4621 
R4 N_11:1 M12:SRC 33.8389 
CC90896 N_11:1 M21:GATE 1.74e-18
CC90928 N_11:1 M5:GATE 2.91e-18
CC90891 N_11:1 A1:1 3.99e-18
CC90917 N_11:1 A2:2 1.691e-17
CC90926 N_11:1 M7:GATE 8.45e-18
CC90925 N_11:1 M6:GATE 7.84e-18
CC90907 N_11:1 M9:GATE 6.03e-18
CC90924 N_11:1 A2 6.219e-17
CC90898 N_11:1 A1 1.082e-17
CC90927 N_11:1 M8:GATE 4.18e-18
CC90899 N_11:1 M12:GATE 3.85e-18
CC90902 N_11:1 M11:GATE 4.99e-18
CC90903 N_11:1 M10:GATE 3.67e-18
CC90966 N_11:1 ZN 9.59e-17
CC90973 N_11:1 M20:SRC 1.14e-18
CC91011 N_11:1 M11:SRC 4.97e-18
CC91019 N_11:1 M9:SRC 4.86e-18
CC90942 N_11:1 ZN:1 1.265e-17
CC90948 N_11:1 ZN:2 8.56e-18
R5 M10:SRC M12:SRC 803.7 
R6 M12:SRC M9:DRN 2001.68 
CC90888 M12:SRC A1:1 3.048e-17
CC90892 M12:SRC A1:2 2.23e-18
CC90913 M12:SRC A2:2 1.21e-18
CC90957 M12:SRC ZN 1.07e-18
R7 M9:DRN M10:SRC 1952.16 
CC90914 M9:DRN A2:2 5.26e-18
CC90906 M9:DRN M9:GATE 2.816e-17
CC90960 M9:DRN ZN 5.69e-18
CC90889 M10:SRC A1:1 7.27e-18
CC90893 M10:SRC A1:2 2.035e-17
CC90904 M10:SRC M10:GATE 9.57e-18
CC90901 M10:SRC M11:GATE 2.999e-17
CC90959 M10:SRC ZN 1.534e-17
CC90916 M5:SRC A2:2 9.26e-18
CC90920 M5:SRC A2:3 6.02e-18
CC90923 M5:SRC A2 1.61e-18
CC90910 M5:SRC A2:1 5.198e-17
CC90912 M5:SRC M20:GATE 5.57e-18
CC90937 M5:SRC ZN:1 3.4e-18
CC90915 M7:SRC A2:2 3.785e-17
CC90911 M7:SRC M20:GATE 5.55e-18
CC90919 M7:SRC A2:3 2.845e-17
CC90922 M7:SRC A2 1.25e-18
C8 N_11:1 0 1.5874e-16
C9 M12:SRC 0 2.27e-17
C10 M9:DRN 0 1.02e-17
C11 M10:SRC 0 8.81e-18
C12 M5:SRC 0 4.4e-18
C13 M7:SRC 0 2.92e-18
R14 A1:1 M23:GATE 266.204 
R15 M11:GATE M23:GATE 1092.88 
R16 M23:GATE A1:2 282.501 
CC91041 M23:GATE N_37:1 6.41e-18
CC91092 M23:GATE M23:SRC 2.937e-17
CC90975 M23:GATE M22:SRC 2.791e-17
CC90950 M23:GATE ZN 1.004e-17
R17 M10:GATE A1:2 94.0755 
R18 M22:GATE A1:2 111.3 
R19 A1:1 A1:2 58.1624 
R20 M11:GATE A1:2 238.78 
R21 M21:GATE A1:2 164.389 
R22 A1:2 M9:GATE 138.947 
CC91017 A1:2 M9:SRC 3.325e-17
CC91010 A1:2 M11:SRC 1.291e-17
CC90964 A1:2 ZN 1.004e-17
R23 M9:GATE M21:GATE 635.948 
CC91108 M21:GATE M21:SRC 2.944e-17
CC91044 M21:GATE N_37:1 6.41e-18
CC90968 M21:GATE M20:SRC 2.802e-17
CC90952 M21:GATE ZN 1.286e-17
R24 M11:GATE A1:1 225.005 
CC90958 M11:GATE ZN 2.77e-18
R25 M12:GATE A1:1 86.5669 
R26 M24:GATE A1:1 111.3 
R27 A1:1 A1 22 
CC91016 A1:1 M9:SRC 1.38e-17
CC91009 A1:1 M11:SRC 3.39e-17
CC91113 A1:1 M21:SRC 1.135e-17
CC91100 A1:1 M23:SRC 1.122e-17
CC91062 A1:1 N_37:1 1.24e-18
CC90963 A1:1 ZN 4.219e-17
CC90986 A1:1 M24:SRC 2.22e-18
CC90980 A1:1 M22:SRC 8.74e-18
CC91008 A1 M11:SRC 1.49e-18
CC91099 A1 M23:SRC 1.82e-18
CC91061 A1 N_37:1 1.04e-18
CC90962 A1 ZN 6.714e-17
CC90985 A1 M24:SRC 2e-18
CC91107 M22:GATE M21:SRC 2.939e-17
CC91043 M22:GATE N_37:1 6.84e-18
CC90976 M22:GATE M22:SRC 2.756e-17
CC90951 M22:GATE ZN 1.275e-17
CC91040 M24:GATE N_37:1 4.03e-18
CC91091 M24:GATE M23:SRC 3e-17
CC90949 M24:GATE ZN 4.74e-18
CC90982 M24:GATE M24:SRC 2.818e-17
CC91006 M12:GATE M11:SRC 2.52e-17
CC91013 M10:GATE M9:SRC 2.505e-17
C28 M23:GATE 0 2.717e-17
C29 A1:2 0 1.68e-17
C30 M9:GATE 0 2.773e-17
C31 M21:GATE 0 4.344e-17
C32 M11:GATE 0 1.987e-17
C33 A1:1 0 1.744e-17
C34 A1 0 1.199e-17
C35 M22:GATE 0 3.087e-17
C36 M24:GATE 0 2.725e-17
C37 M12:GATE 0 1.713e-17
C38 M10:GATE 0 2.291e-17
R39 M17:GATE A2:1 111.3 
CC91132 M17:GATE M17:SRC 9.37e-18
CC91050 M17:GATE N_37:1 6.06e-18
CC90956 M17:GATE ZN 3.02e-18
CC90999 M17:GATE M17:DRN 4.87e-18
CC90934 M17:GATE ZN:1 1.95e-18
R40 A2 A2:1 22.4117 
R41 M5:GATE A2:1 110.162 
R42 M6:GATE A2:1 141.186 
R43 A2:1 A2:3 29.4771 
CC91139 A2:1 M17:SRC 2.004e-17
CC91004 A2:1 M17:DRN 2.342e-17
R44 A2 A2:3 22.2732 
R45 M6:GATE A2:3 340.795 
R46 M7:GATE A2:3 82.8124 
R47 A2:2 A2:3 24.9722 
R48 A2:3 M18:GATE 111.3 
CC91049 M18:GATE N_37:1 6.74e-18
CC90955 M18:GATE ZN 3.75e-18
CC91131 M18:GATE M17:SRC 2.948e-17
CC90990 M18:GATE M18:SRC 2.814e-17
CC90933 M18:GATE ZN:1 1.05e-18
R49 M19:GATE A2:2 111.3 
R50 A2 A2:2 22.1375 
R51 M8:GATE A2:2 86.5669 
R52 A2:2 M20:GATE 133.466 
CC90972 A2:2 M20:SRC 2.84e-17
CC91138 A2:2 M17:SRC 4.6e-18
CC90947 A2:2 ZN:2 1.469e-17
CC91126 A2:2 M19:SRC 4.51e-17
CC90965 A2:2 ZN 3.47e-18
CC90994 A2:2 M18:SRC 5.81e-18
CC91102 A2:2 M23:SRC 1.114e-17
CC91003 A2:2 M17:DRN 4.89e-18
CC90988 M20:GATE M18:SRC 4.25e-18
CC91128 M20:GATE M17:SRC 8.08e-18
CC91119 M20:GATE M19:SRC 1.724e-17
CC91046 M20:GATE N_37:1 1.41e-18
CC90997 M20:GATE M17:DRN 2.86e-18
CC90932 M20:GATE ZN:1 4.36e-18
CC90938 M5:GATE ZN:1 3.57e-18
CC91060 A2 N_37:1 4.01e-18
CC90961 A2 ZN 4.064e-17
CC91002 A2 M17:DRN 1.27e-18
CC90939 A2 ZN:1 1.965e-17
CC90989 M19:GATE M18:SRC 2.808e-17
CC91047 M19:GATE N_37:1 1.46e-18
CC91120 M19:GATE M19:SRC 9.46e-18
C53 M17:GATE 0 2.801e-17
C54 A2:1 0 1.584e-17
C55 A2:3 0 1.528e-17
C56 M18:GATE 0 3.482e-17
C57 A2:2 0 5.288e-17
C58 M20:GATE 0 4.148e-17
C59 M8:GATE 0 3.678e-17
C60 M7:GATE 0 3.223e-17
C61 M6:GATE 0 4.197e-17
C62 M5:GATE 0 5.547e-17
C63 A2 0 2.228e-17
C64 M19:GATE 0 2.307e-17
R65 M12:DRN M11:SRC 0.001 
R66 M11:SRC ZN 30.3374 
R67 M24:SRC ZN 40.0778 
R68 M9:SRC ZN 30.3702 
R69 ZN:2 ZN 0.92654 
R70 ZN M22:SRC 39.0574 
CC91058 ZN N_37:1 1.7741e-16
CC91135 ZN M17:SRC 4.5e-18
CC91123 ZN M19:SRC 4.5e-18
CC91112 ZN M21:SRC 5.39e-18
CC91098 ZN M23:SRC 4.67e-18
R71 M23:DRN M22:SRC 0.001 
R72 M22:SRC ZN:2 135.425 
CC91042 M22:SRC N_37:1 6.6e-18
R73 M20:SRC ZN:2 29.9999 
R74 M24:SRC ZN:2 135.741 
R75 M18:SRC ZN:2 41.1421 
R76 ZN:1 ZN:2 2.95584 
R77 ZN:2 M17:DRN 66.1317 
CC91063 ZN:2 N_37:1 4.715e-17
CC91101 ZN:2 M23:SRC 7.45e-18
CC91125 ZN:2 M19:SRC 1.249e-17
CC91114 ZN:2 M21:SRC 1.945e-17
CC91029 ZN:2 B 6.5e-18
CC91022 ZN:2 B:1 8.14e-18
R78 M17:DRN ZN:1 58.5751 
CC91034 M17:DRN M16:GATE 3.57e-18
CC91051 M17:DRN N_37:1 7.34e-18
R79 M1:SRC ZN:1 30.5689 
R80 M3:SRC ZN:1 29.9999 
R81 ZN:1 M18:SRC 118.609 
CC91065 ZN:1 N_37:1 1.171e-17
CC91038 ZN:1 M4:GATE 4.57e-18
CC91036 ZN:1 M16:GATE 1.303e-17
CC91103 ZN:1 M23:SRC 1.32e-18
CC91078 ZN:1 M15:SRC 1.3e-18
CC91031 ZN:1 M2:GATE 8.1e-18
CC91030 ZN:1 B 6.366e-17
CC91032 ZN:1 M1:GATE 2.02e-18
R82 M18:SRC M19:DRN 0.001 
CC91048 M18:SRC N_37:1 6.6e-18
R83 M9:SRC M10:DRN 0.001 
R84 M20:SRC M21:DRN 0.001 
CC91045 M20:SRC N_37:1 6.6e-18
R85 M3:SRC M4:DRN 0.001 
CC91037 M3:SRC M4:GATE 2.412e-17
CC91033 M3:SRC M3:GATE 8.65e-18
CC91027 M3:SRC B 1.946e-17
CC91020 M3:SRC B:1 1.99e-17
R86 M1:SRC M2:DRN 0.001 
CC91025 M1:SRC B:2 2.854e-17
CC91028 M1:SRC B 4.401e-17
C87 M11:SRC 0 2.48e-18
C88 ZN 0 3.017e-17
C89 M22:SRC 0 4.03e-18
C90 ZN:2 0 1.739e-17
C91 M17:DRN 0 1.817e-17
C92 ZN:1 0 7.391e-17
C93 M18:SRC 0 3.26e-18
C94 M9:SRC 0 7.35e-18
C95 M24:SRC 0 2.476e-17
C96 M20:SRC 0 1.87e-18
C97 M3:SRC 0 8.28e-18
C98 M1:SRC 0 2.96e-18
R99 M2:GATE B:2 94.0755 
R100 M14:GATE B:2 111.3 
R101 B:1 B:2 27.6389 
R102 B B:2 23.3574 
R103 M13:GATE B:2 259.177 
R104 B:2 M1:GATE 187.595 
CC91089 B:2 M13:SRC 1.082e-17
R105 B M1:GATE 208.822 
R106 M1:GATE M13:GATE 1038.31 
R107 M13:GATE B 288.505 
CC91055 M13:GATE N_37:1 5.29e-18
CC91084 M13:GATE M13:SRC 4.421e-17
R108 M4:GATE B 529.497 
R109 M16:GATE B 499.665 
R110 B B:1 23.0871 
CC91087 B M13:SRC 1.64e-18
CC91059 B N_37:1 5.081e-17
CC91076 B M15:SRC 1.29e-18
R111 M15:GATE B:1 111.3 
R112 M3:GATE B:1 94.0755 
R113 M4:GATE B:1 190.021 
R114 B:1 M16:GATE 179.317 
CC91088 B:1 M13:SRC 9.67e-18
CC91079 B:1 M15:SRC 1.876e-17
R115 M16:GATE M4:GATE 558.737 
CC91070 M16:GATE M15:SRC 4.655e-17
CC91052 M16:GATE N_37:1 1.181e-17
CC91056 M4:GATE N_37:1 1.71e-18
CC91073 M4:GATE M15:SRC 4.46e-18
CC91085 M4:GATE M13:SRC 4.35e-18
CC91095 M15:GATE M23:SRC 5.95e-18
CC91071 M15:GATE M15:SRC 4.548e-17
CC91053 M15:GATE N_37:1 4.9e-18
CC91096 M14:GATE M23:SRC 2.37e-18
CC91054 M14:GATE N_37:1 8.01e-18
CC91083 M14:GATE M13:SRC 4.53e-17
C116 M2:GATE 0 3.544e-17
C117 B:2 0 2.488e-17
C118 M1:GATE 0 5.74e-17
C119 M13:GATE 0 7.77e-17
C120 B 0 3.705e-17
C121 B:1 0 5.556e-17
C122 M16:GATE 0 6.335e-17
C123 M4:GATE 0 4.782e-17
C124 M3:GATE 0 3.315e-17
C125 M15:GATE 0 2.909e-17
C126 M14:GATE 0 3.457e-17
R127 N_37:1 M23:SRC 34.4635 
R128 M19:SRC M23:SRC 1418.07 
R129 M23:SRC M21:SRC 700.523 
R130 N_37:1 M21:SRC 33.6459 
R131 M21:SRC M19:SRC 1384.42 
R132 M19:SRC N_37:1 32.1037 
R133 M13:SRC N_37:1 17.993 
R134 M15:SRC N_37:1 17.109 
R135 N_37:1 M17:SRC 29.9999 
R136 M15:SRC M13:SRC 267.739 
C137 M23:SRC 0 1.512e-17
C138 M21:SRC 0 1.727e-17
C139 M19:SRC 0 5.86e-18
C140 N_37:1 0 2.5562e-16
C141 M17:SRC 0 5.86e-18
C142 M15:SRC 0 2.41e-17
C143 M13:SRC 0 1.567e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
