.SUBCKT OR2D1 A1 A2 Z
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.8e-14  AS=5.8e-14  PD=1.13e-06  PS=8.53e-07  SA=3.28e-07  SB=1.75e-07  NRD=0.496  NRS=0.755  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=2.04e-07  AD=2.9e-14  AS=2e-14  PD=4.27e-07  PS=4.05e-07  SA=4.7e-07  SB=4.85e-07  NRD=0.882  NRS=5.196  SCA=18.109  SCB=0.02  SCC=0.002 
MMM3 M2:SRC M3:GATE vss vss nch L=6e-08 W=2.04e-07  AD=2e-14  AS=3.9e-14  PD=4.05e-07  PS=7.9e-07  SA=2e-07  SB=7.55e-07  NRD=5.196  NRS=1.534  SCA=18.109  SCB=0.02  SCC=0.002 
MMM4 M4:DRN M4:GATE vdd vdd pch L=6e-08 W=5.23e-07  AD=9.1e-14  AS=7.3e-14  PD=1.39e-06  PS=8e-07  SA=7.75e-07  SB=1.75e-07  NRD=0.446  NRS=0.644  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=5.24e-07  AD=7.3e-14  AS=5.2e-14  PD=8e-07  PS=7.2e-07  SA=4.35e-07  SB=5.15e-07  NRD=0.644  NRS=2.009  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M5:SRC M6:GATE M6:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=9.1e-14  PD=7.2e-07  PS=1.39e-06  SA=1.75e-07  SB=7.75e-07  NRD=2.009  NRS=0.446  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M4:DRN Z 15.4724 
R1 Z M1:DRN 15.266 
CC10664 Z M4:GATE 5.52e-18
CC10667 Z M6:SRC 8.23e-17
CC10669 Z M1:GATE 1.027e-17
CC10666 M1:DRN M6:SRC 4.086e-17
CC10668 M1:DRN M1:GATE 9.66e-18
CC10665 M4:DRN M6:SRC 1.65e-18
CC10663 M4:DRN M4:GATE 4.785e-17
C2 Z 0 1.0224e-16
C3 M1:DRN 0 2.251e-17
C4 M4:DRN 0 3.155e-17
R5 M4:GATE M2:SRC 488.309 
R6 M6:SRC M2:SRC 54.8362 
R7 M2:SRC M1:GATE 401.352 
CC10678 M2:SRC M2:GATE 9.16e-18
CC10691 M2:SRC M3:GATE 1.158e-17
CC10686 M2:SRC A1 3.449e-17
CC10675 M2:SRC A2 1.2517e-16
R8 M4:GATE M1:GATE 411.537 
R9 M1:GATE M6:SRC 212.732 
CC10679 M1:GATE M2:GATE 1.97e-18
CC10688 M1:GATE A1 1.469e-17
CC10676 M1:GATE A2 2.13e-18
R10 M6:SRC M4:GATE 258.825 
CC10680 M6:SRC M6:GATE 5.591e-17
CC10677 M6:SRC M2:GATE 1.25e-17
CC10690 M6:SRC M3:GATE 6.16e-18
CC10684 M6:SRC A1 2.182e-17
CC10671 M6:SRC M5:GATE 1.245e-17
CC10674 M4:GATE A2 1.152e-17
CC10672 M4:GATE M5:GATE 4.32e-18
C11 M2:SRC 0 3.214e-17
C12 M1:GATE 0 7.416e-17
C13 M6:SRC 0 1.2063e-16
C14 M4:GATE 0 9.682e-17
R15 M5:GATE M2:GATE 385.604 
R16 M2:GATE A2 87.7049 
CC10692 M2:GATE M3:GATE 1.86e-18
CC10687 M2:GATE A1 1.57e-18
R17 A2 M5:GATE 158.476 
CC10693 A2 M3:GATE 4.83e-18
CC10683 A2 M6:GATE 3.8e-18
CC10689 A2 A1 2.911e-17
CC10685 M5:GATE A1 1.129e-17
CC10681 M5:GATE M6:GATE 1.374e-17
C18 M2:GATE 0 3.27e-17
C19 A2 0 8.83e-18
C20 M5:GATE 0 7.494e-17
R21 M3:GATE A1 86.6423 
R22 A1 M6:GATE 158.15 
R23 M6:GATE M3:GATE 373.471 
C24 A1 0 5.084e-17
C25 M6:GATE 0 4.944e-17
C26 M3:GATE 0 2.947e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
