.SUBCKT ND2D8 A1 A2 ZN
MMM20 M20:DRN M20:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.26e-06  SB=9.4e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 vdd M21:GATE M21:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3e-06  SB=1.2e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.74e-06  SB=1.46e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 vdd M23:GATE M23:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.48e-06  SB=1.72e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 vdd M24:GATE M24:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.72e-06  SB=2.48e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM25 vdd M25:GATE M25:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.46e-06  SB=2.74e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM26 M26:DRN M26:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=2.22e-06  SB=1.98e-06  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM27 M27:DRN M27:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.98e-06  SB=2.22e-06  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM28 M28:DRN M28:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.2e-06  SB=3e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM29 vdd M29:GATE M29:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.4e-07  SB=3.26e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M7:SRC M10:GATE vss vss nch L=6e-08 W=2.3e-07  AD=2.3e-14  AS=2.3e-14  PD=4.3e-07  PS=4.3e-07  SA=2.24e-06  SB=1.96e-06  NRD=6.986  NRS=7.015  SCA=16.543  SCB=0.019  SCC=0.002 
MMM11 M9:SRC M11:GATE vss vss nch L=6e-08 W=2.3e-07  AD=2.3e-14  AS=2.3e-14  PD=4.3e-07  PS=4.3e-07  SA=1.98e-06  SB=2.22e-06  NRD=6.986  NRS=7.015  SCA=16.543  SCB=0.019  SCC=0.002 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=8e-14  AS=4.4e-14  PD=1.19e-06  PS=6.15e-07  SA=2.261e-06  SB=2.05e-07  NRD=0.566  NRS=0.288  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M8:SRC M12:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.2e-06  SB=8.57e-07  NRD=4.12  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M1:SRC M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=4.4e-14  AS=3.9e-14  PD=6.15e-07  PS=5.9e-07  SA=1.89e-06  SB=4.9e-07  NRD=0.288  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.4e-07  SB=1.277e-06  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.53e-06  SB=7.5e-07  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M13:SRC M14:GATE M14:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=1.655e-06  NRD=4.12  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M3:SRC M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=1.139e-06  SB=1.01e-06  NRD=4.12  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 M15:DRN M15:GATE M15:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=2.006e-06  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=2.5e-14  PD=5.7e-07  PS=5.2e-07  SA=7.35e-07  SB=1.25e-06  NRD=7.648  NRS=14.848  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 vss M16:GATE M15:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.6e-07  SB=2.339e-06  NRD=0.462  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M5:SRC M6:GATE M6:SRC vss nch L=6e-08 W=3.9e-07  AD=2.5e-14  AS=4.4e-14  PD=5.2e-07  PS=7.42e-07  SA=3.72e-07  SB=1.44e-06  NRD=14.848  NRS=7.393  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 vdd M17:GATE M17:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=4.04e-06  SB=1.6e-07  NRD=0.427  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 M7:DRN M7:GATE M7:SRC vss nch L=6e-08 W=2.36e-07  AD=2.6e-14  AS=2.3e-14  PD=4.38e-07  PS=4.3e-07  SA=2.5e-06  SB=1.7e-06  NRD=0.51  NRS=6.986  SCA=16.543  SCB=0.019  SCC=0.002 
MMM18 M18:DRN M18:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.78e-06  SB=4.2e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE M8:SRC vss nch L=6e-08 W=3.9e-07  AD=4.4e-14  AS=3.9e-14  PD=7.42e-07  PS=5.9e-07  SA=1.46e-06  SB=3.71e-07  NRD=7.393  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vdd M19:GATE M19:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.52e-06  SB=6.8e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 M9:DRN M9:GATE M9:SRC vss nch L=6e-08 W=2.36e-07  AD=2.6e-14  AS=2.3e-14  PD=4.38e-07  PS=4.3e-07  SA=1.72e-06  SB=2.48e-06  NRD=0.51  NRS=6.986  SCA=16.543  SCB=0.019  SCC=0.002 
MMM30 M30:DRN M30:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=3.52e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM31 vdd M31:GATE M31:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=3.78e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM32 M32:DRN M32:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=4.04e-06  NRD=2.099  NRS=0.427  SCA=9.643  SCB=0.01  SCC=0.000823 
CC45318 M1:SRC A1:2 2.05e-18
CC45203 M3:SRC A2:1 2.07e-18
CC45457 M7:SRC M7:GATE 1.47e-18
CC45454 M9:SRC M7:GATE 1.47e-18
R0 M22:DRN M21:SRC 0.001 
R1 ZN:4 M21:SRC 61.1029 
R2 M21:SRC ZN:2 60.3402 
CC45308 M21:SRC A1:2 6.56e-18
CC45349 M21:SRC M22:GATE 2.784e-17
CC45236 M21:SRC M21:GATE 2.823e-17
CC45200 M21:SRC A2:1 3.21e-18
R3 M7:DRN ZN:2 194.098 
R4 M17:SRC ZN:2 31.2033 
R5 M19:SRC ZN:2 29.9999 
R6 ZN:4 ZN:2 1.46695 
R7 ZN:2 M2:SRC 32.2118 
CC45385 ZN:2 M3:GATE 2.44e-18
CC45304 ZN:2 A1:1 5.818e-17
CC45378 ZN:2 M2:GATE 6.29e-18
CC45322 ZN:2 A1:2 1.486e-17
CC45368 ZN:2 M18:GATE 1.998e-17
CC45362 ZN:2 M19:GATE 2.91e-18
CC45226 ZN:2 A2:4 7.47e-18
CC45233 ZN:2 A2:5 1.194e-17
CC45238 ZN:2 M21:GATE 1.04e-18
CC45244 ZN:2 M17:GATE 3.96e-18
CC45252 ZN:2 M32:GATE 1.141e-17
CC45214 ZN:2 A2:2 6.233e-17
R8 M17:SRC M2:SRC 1952.36 
R9 M2:SRC M3:DRN 0.001 
CC45383 M2:SRC M3:GATE 1.48e-18
CC45317 M2:SRC A1:2 7.358e-17
CC45212 M2:SRC A2:2 9.99e-18
R10 M9:DRN ZN:1 31.1786 
R11 M29:SRC ZN:1 96.7371 
R12 M25:SRC ZN:1 42.4842 
R13 M27:DRN ZN:1 48.6908 
R14 ZN ZN:1 0.54731 
R15 ZN:1 ZN:3 1.85348 
CC45413 ZN:1 M25:GATE 1.14e-18
CC45227 ZN:1 A2:4 1.54e-18
CC45234 ZN:1 A2:5 1.15e-18
CC45423 ZN:1 M24:GATE 6.78e-18
CC45215 ZN:1 A2:2 7.02e-18
CC45270 ZN:1 M27:GATE 1.29e-18
CC45490 ZN:1 M9:GATE 1.521e-17
CC45479 ZN:1 M8:GATE 1.9e-18
CC45284 ZN:1 A2 8.261e-17
CC45445 ZN:1 A1 4.638e-17
R16 M29:SRC ZN:3 44.3122 
R17 M31:SRC ZN:3 30.1454 
R18 M25:SRC ZN:3 108.502 
R19 ZN:3 M14:SRC 31.236 
CC45333 ZN:3 A1:3 9.65e-18
CC45404 ZN:3 M30:GATE 2.79e-18
CC45216 ZN:3 A2:2 2.705e-17
CC45394 ZN:3 M31:GATE 5.62e-18
CC45253 ZN:3 M32:GATE 9.48e-18
CC45475 ZN:3 M15:GATE 5.88e-18
CC45287 ZN:3 M16:GATE 1.31e-18
CC45285 ZN:3 A2 5.583e-17
CC45446 ZN:3 A1 5.219e-17
R20 M14:SRC M15:DRN 0.001 
CC45330 M14:SRC A1:3 6.37e-17
CC45439 M14:SRC A1 1.22e-17
CC45282 M14:SRC A2 8.57e-18
R21 M7:DRN ZN:4 37.5642 
R22 M23:SRC ZN:4 29.9999 
R23 ZN:4 ZN 0.05576 
CC45373 ZN:4 M6:GATE 3.12e-18
CC45306 ZN:4 A1:1 2.768e-17
CC45379 ZN:4 M2:GATE 5.24e-18
CC45334 ZN:4 A1:3 1.63e-18
CC45354 ZN:4 M22:GATE 4.67e-18
CC45324 ZN:4 A1:2 1.0063e-16
CC45363 ZN:4 M19:GATE 4.32e-18
CC45260 ZN:4 M29:GATE 4.77e-18
CC45235 ZN:4 A2:5 2.09e-18
CC45405 ZN:4 M30:GATE 4.13e-18
CC45239 ZN:4 M21:GATE 3.9e-18
CC45425 ZN:4 M24:GATE 3.78e-18
CC45271 ZN:4 M27:GATE 3.47e-18
CC45217 ZN:4 A2:2 2.097e-17
CC45223 ZN:4 A2:3 1.5e-18
CC45415 ZN:4 M25:GATE 4.14e-18
CC45265 ZN:4 M28:GATE 4.14e-18
CC45395 ZN:4 M31:GATE 4.1e-18
CC45242 ZN:4 M20:GATE 4.1e-18
CC45254 ZN:4 M32:GATE 2.38e-18
CC45245 ZN:4 M17:GATE 2.38e-18
CC45464 ZN:4 M7:GATE 1.508e-17
CC45491 ZN:4 M9:GATE 1.8e-18
CC45277 ZN:4 M26:GATE 3.35e-18
CC45434 ZN:4 M23:GATE 1.185e-17
CC45286 ZN:4 A2 8.045e-17
CC45447 ZN:4 A1 1.0786e-16
CC45205 ZN:4 A2:1 1.52e-18
R24 ZN M27:DRN 79.0308 
CC45232 ZN A2:5 5.35e-18
CC45268 ZN M27:GATE 4.2e-18
CC45432 ZN M23:GATE 1.48e-18
CC45274 ZN M26:GATE 8.53e-18
CC45213 ZN A2:2 2.277e-17
R25 M27:DRN M24:SRC 0.001 
CC45418 M27:DRN M24:GATE 2.815e-17
CC45266 M27:DRN M27:GATE 2.821e-17
CC45206 M27:DRN A2:2 1.68e-18
R26 M19:SRC M20:DRN 0.001 
CC45375 M19:SRC M2:GATE 1.68e-18
CC45311 M19:SRC A1:2 2.85e-18
CC45358 M19:SRC M19:GATE 2.765e-17
CC45240 M19:SRC M20:GATE 8.15e-18
CC45294 M19:SRC A1:1 6.42e-18
CC45208 M19:SRC A2:2 2.016e-17
R27 M17:SRC M18:DRN 0.001 
CC45366 M17:SRC M18:GATE 2.8e-17
CC45243 M17:SRC M17:GATE 2.839e-17
CC45249 M17:SRC M1:GATE 1.11e-18
CC45209 M17:SRC A2:2 3.08e-18
R28 M28:DRN M25:SRC 0.001 
CC45262 M25:SRC M28:GATE 2.821e-17
CC45410 M25:SRC M25:GATE 2.789e-17
CC45438 M25:SRC A1 6.53e-18
R29 M26:DRN M23:SRC 0.001 
CC45230 M23:SRC A2:5 1.53e-18
CC45429 M23:SRC M23:GATE 2.789e-17
CC45281 M23:SRC A2 1.5e-18
CC45273 M23:SRC M26:GATE 2.76e-17
R30 M31:SRC M32:DRN 0.001 
CC45388 M31:SRC M31:GATE 2.785e-17
CC45251 M31:SRC M32:GATE 2.835e-17
CC45278 M31:SRC A2 1.03e-18
R31 M6:SRC M7:DRN 0.001 
CC45314 M7:DRN A1:2 1.09e-18
CC45458 M7:DRN M7:GATE 2.477e-17
CC45297 M7:DRN A1:1 4.938e-17
CC45485 M7:DRN M9:GATE 6.78e-18
CC45290 M7:DRN M10:GATE 1.64e-18
CC45211 M7:DRN A2:2 4.23e-18
R32 M29:SRC M30:DRN 0.001 
CC45255 M29:SRC M29:GATE 2.766e-17
CC45398 M29:SRC M30:GATE 2.803e-17
CC45435 M29:SRC A1 6.17e-18
CC45279 M29:SRC A2 1.09e-18
R33 M8:DRN M9:DRN 0.001 
CC45339 M9:DRN A1:4 5.104e-17
CC45289 M9:DRN M11:GATE 1.64e-18
CC45484 M9:DRN M9:GATE 3.135e-17
CC45283 M9:DRN A2 6.39e-18
CC45440 M9:DRN A1 1.24e-18
C34 M21:SRC 0 9.23e-18
C35 ZN:2 0 7.46e-18
C36 M2:SRC 0 4.47e-18
C37 ZN:1 0 8.24e-18
C38 ZN:3 0 1.438e-17
C39 M14:SRC 0 3.4e-18
C40 ZN:4 0 4.0252e-16
C41 ZN 0 3.38e-17
C42 M27:DRN 0 3.92e-18
C43 M19:SRC 0 1.569e-17
C44 M17:SRC 0 1.677e-17
C45 M25:SRC 0 8.83e-18
C46 M23:SRC 0 4e-18
C47 M31:SRC 0 5.82e-18
C48 M7:DRN 0 1.52e-17
C49 M29:SRC 0 8.65e-18
C50 M9:DRN 0 1.524e-17
R51 A2:2 M32:GATE 1977.64 
R52 A2 M32:GATE 163.037 
R53 M32:GATE M16:GATE 462.455 
CC45387 M32:GATE M31:GATE 7.97e-18
R54 A2:2 M16:GATE 1617.57 
R55 M16:GATE A2 133.352 
CC45472 M16:GATE M15:GATE 4.15e-18
CC45329 M16:GATE A1:3 1.165e-17
R56 M12:GATE A2 220.204 
R57 M28:GATE A2 300.988 
R58 A2:2 A2 5.13701 
R59 A2:3 A2 48.1172 
R60 A2:5 A2 102.494 
R61 A2 A2:4 166.551 
CC45460 A2 M7:GATE 4.57e-18
CC45442 A2 A1 6.431e-17
CC45487 A2 M9:GATE 6.27e-18
CC45478 A2 M8:GATE 2.29e-18
CC45474 A2 M15:GATE 9.53e-18
CC45469 A2 M14:GATE 7.98e-18
CC45401 A2 M30:GATE 1.91e-18
CC45341 A2 A1:4 1.186e-17
CC45331 A2 A1:3 8.86e-18
CC45300 A2 A1:1 3.85e-18
R62 M11:GATE A2:4 72.8752 
R63 M27:GATE A2:4 111.3 
R64 A2:2 A2:4 122.949 
R65 A2:4 A2:5 18.4701 
CC45488 A2:4 M9:GATE 1.82e-18
CC45343 A2:4 A1:4 1.87e-18
R66 M10:GATE A2:5 72.8752 
R67 A2:2 A2:5 75.6607 
R68 A2:5 M26:GATE 111.3 
CC45461 A2:5 M7:GATE 2.42e-18
CC45344 A2:5 A1:4 7.68e-18
CC45302 A2:5 A1:1 9.5e-18
CC45428 M26:GATE M23:GATE 7.71e-18
R69 M13:GATE A2:3 94.0755 
R70 M12:GATE A2:3 178.093 
R71 M28:GATE A2:3 243.428 
R72 A2:3 M29:GATE 111.3 
CC45443 A2:3 A1 9.56e-18
CC45470 A2:3 M14:GATE 4.29e-18
CC45411 A2:3 M25:GATE 1.32e-18
CC45342 A2:3 A1:4 7.59e-18
CC45332 A2:3 A1:3 8.25e-18
CC45436 M29:GATE A1 4.22e-18
CC45399 M29:GATE M30:GATE 7.53e-18
CC45328 M29:GATE A1:3 1.26e-18
R73 M5:GATE A2:1 92.75 
CC45370 M5:GATE M6:GATE 6.39e-18
CC45298 M5:GATE A1:1 8.17e-18
R74 A2:2 A2:1 50.3476 
R75 M20:GATE A2:1 252.457 
R76 M4:GATE A2:1 192.065 
R77 A2:1 M21:GATE 112.625 
CC45462 A2:1 M7:GATE 7.56e-18
CC45321 A2:1 A1:2 1.886e-17
CC45372 A2:1 M6:GATE 6.02e-18
CC45303 A2:1 A1:1 9.59e-18
CC45350 M21:GATE M22:GATE 7.66e-18
CC45309 M21:GATE A1:2 4.96e-18
R78 A2:2 M4:GATE 226.097 
R79 M4:GATE M20:GATE 1133.71 
CC45382 M4:GATE M3:GATE 3.84e-18
CC45316 M4:GATE A1:2 9.26e-18
CC45299 M4:GATE A1:1 2.39e-18
R80 M20:GATE A2:2 297.19 
CC45357 M20:GATE M19:GATE 7.25e-18
CC45310 M20:GATE A1:2 3.33e-18
CC45293 M20:GATE A1:1 5.42e-18
R81 M1:GATE A2:2 124.045 
R82 A2:2 M17:GATE 150.568 
CC45465 A2:2 M7:GATE 3.56e-18
CC45448 A2:2 A1 7.49e-18
CC45426 A2:2 M24:GATE 3.35e-18
CC45492 A2:2 M9:GATE 1.353e-17
CC45480 A2:2 M8:GATE 5.85e-18
CC45325 A2:2 A1:2 1.13e-17
CC45386 A2:2 M3:GATE 9.72e-18
CC45380 A2:2 M2:GATE 2.02e-17
CC45374 A2:2 M6:GATE 7.97e-18
CC45307 A2:2 A1:1 5.401e-17
R83 M17:GATE M1:GATE 508.741 
CC45367 M17:GATE M18:GATE 3.77e-18
CC45313 M17:GATE A1:2 4.18e-18
CC45377 M1:GATE M2:GATE 3.69e-18
CC45319 M1:GATE A1:2 1.249e-17
CC45417 M27:GATE M24:GATE 7.89e-18
R84 M28:GATE M12:GATE 1114.02 
CC45437 M28:GATE A1 5.28e-18
CC45407 M28:GATE M25:GATE 7.78e-18
CC45477 M12:GATE M8:GATE 4.16e-18
CC45337 M12:GATE A1:4 8.21e-18
CC45455 M10:GATE M7:GATE 1.136e-17
CC45453 M11:GATE M7:GATE 3.17e-18
CC45482 M11:GATE M9:GATE 8.4e-18
CC45467 M13:GATE M14:GATE 7.75e-18
C85 M32:GATE 0 8.183e-17
C86 M16:GATE 0 5.034e-17
C87 A2 0 3.3173e-16
C88 A2:4 0 2.047e-17
C89 A2:5 0 5.373e-17
C90 M26:GATE 0 5.161e-17
C91 A2:3 0 5.476e-17
C92 M29:GATE 0 6.761e-17
C93 M5:GATE 0 2.039e-17
C94 A2:1 0 5.553e-17
C95 M21:GATE 0 4.678e-17
C96 M4:GATE 0 2.05e-17
C97 M20:GATE 0 3.313e-17
C98 A2:2 0 3.3413e-16
C99 M17:GATE 0 8.545e-17
C100 M1:GATE 0 3.322e-17
C101 M27:GATE 0 4.893e-17
C102 M28:GATE 0 6.17e-17
C103 M12:GATE 0 2.926e-17
C104 M10:GATE 0 2.681e-17
C105 M11:GATE 0 2.692e-17
C106 M13:GATE 0 4.274e-17
R107 M19:GATE A1:2 111.3 
R108 M3:GATE A1:2 80.5597 
R109 A1:1 A1:2 45.7303 
R110 M2:GATE A1:2 130.628 
R111 A1:2 M18:GATE 159.74 
R112 M18:GATE M2:GATE 747.315 
R113 M22:GATE A1:1 111.3 
R114 M6:GATE A1:1 83.8364 
R115 M7:GATE A1:1 84.1834 
R116 A1:1 M23:GATE 176.674 
R117 M23:GATE M7:GATE 388.204 
R118 M7:GATE M9:GATE 413.402 
R119 M24:GATE M9:GATE 438.154 
R120 M9:GATE A1:4 70.0443 
R121 M8:GATE A1:4 81.4271 
R122 M24:GATE A1:4 173.052 
R123 A1 A1:4 23.8381 
R124 A1:4 M25:GATE 111.3 
R125 M15:GATE A1:3 94.0755 
R126 M31:GATE A1:3 111.3 
R127 M14:GATE A1:3 162.232 
R128 M30:GATE A1:3 233.348 
R129 A1:3 A1 46.1243 
R130 M14:GATE A1 219.252 
R131 A1 M30:GATE 315.362 
R132 M30:GATE M14:GATE 1109.22 
C133 M19:GATE 0 5.902e-17
C134 A1:2 0 3.416e-17
C135 M18:GATE 0 2.678e-17
C136 M2:GATE 0 3.921e-17
C137 M22:GATE 0 5.125e-17
C138 A1:1 0 1.829e-17
C139 M23:GATE 0 8.467e-17
C140 M7:GATE 0 1.1506e-16
C141 M9:GATE 0 3.841e-17
C142 A1:4 0 1.308e-17
C143 M25:GATE 0 6.808e-17
C144 A1:3 0 1.887e-17
C145 A1 0 1.266e-17
C146 M30:GATE 0 6.942e-17
C147 M14:GATE 0 2.675e-17
C148 M24:GATE 0 8.223e-17
C149 M31:GATE 0 6.609e-17
C150 M3:GATE 0 2.076e-17
C151 M6:GATE 0 2.057e-17
C152 M15:GATE 0 2.638e-17
C153 M8:GATE 0 2.767e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
