.SUBCKT XOR2D2 A1 A2 Z
MMM10 vdd M10:GATE M10:SRC vdd pch L=6e-08 W=2.64e-07  AD=4.5e-14  AS=4.2e-14  PD=7.45e-07  PS=8.4e-07  SA=1.6e-07  SB=1.75e-07  NRD=0.684  NRS=0.704  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=9.23e-07  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.081e-06  SB=1.6e-07  NRD=0.567  NRS=4.141  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.8e-14  PD=7.2e-07  PS=7.45e-07  SA=6.4e-07  SB=4.2e-07  NRD=2.099  NRS=0.296  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.81e-07  SB=4.2e-07  NRD=4.141  NRS=4.183  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.21e-07  AD=5.8e-14  AS=7.1e-14  PD=7.45e-07  PS=9.49e-07  SA=3.08e-07  SB=7.05e-07  NRD=0.296  NRS=0.341  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4.1e-14  PD=5.9e-07  PS=6.48e-07  SA=4.25e-07  SB=6.8e-07  NRD=4.183  NRS=5.861  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM14 M8:SRC M14:GATE M13:SRC vdd pch L=6e-08 W=3.47e-07  AD=4.9e-14  AS=4.6e-14  PD=8e-07  PS=6.21e-07  SA=1.96e-07  SB=8.04e-07  NRD=0.459  NRS=0.43  SCA=4.486  SCB=0.003  SCC=4.492e-05 
MMM4 M3:SRC M4:GATE M4:SRC vss nch L=6e-08 W=3.28e-07  AD=3.3e-14  AS=4.3e-14  PD=5.32e-07  PS=6.45e-07  SA=3.73e-07  SB=9.4e-07  NRD=0.366  NRS=0.46  SCA=11.685  SCB=0.013  SCC=0.000978 
MMM5 M4:SRC M5:GATE M5:SRC vss nch L=6e-08 W=3.19e-07  AD=4.2e-14  AS=4.6e-14  PD=6.25e-07  PS=8.43e-07  SA=1.78e-07  SB=5.64e-07  NRD=0.471  NRS=0.521  SCA=7.393  SCB=0.008  SCC=0.0002747 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=1.99e-07  AD=3.5e-14  AS=2.1e-14  PD=7.5e-07  PS=4.25e-07  SA=1.8e-07  SB=4.79e-07  NRD=0.972  NRS=5.674  SCA=14.747  SCB=0.017  SCC=0.001 
MMM7 M5:SRC M7:GATE vss vss nch L=6.2e-08 W=1.93e-07  AD=2.8e-14  AS=2e-14  PD=5.17e-07  PS=4.15e-07  SA=3.58e-07  SB=3.87e-07  NRD=0.799  NRS=4.081  SCA=18.359  SCB=0.02  SCC=0.002 
MMM8 M8:DRN M8:GATE M8:SRC vdd pch L=6e-08 W=3.13e-07  AD=3.2e-14  AS=4.4e-14  PD=5.55e-07  PS=7.3e-07  SA=3.23e-07  SB=2.63e-07  NRD=7.25  NRS=0.493  SCA=13.685  SCB=0.015  SCC=0.001 
MMM9 M8:DRN M9:GATE vdd vdd pch L=6e-08 W=2.66e-07  AD=2.7e-14  AS=4.5e-14  PD=4.65e-07  PS=7.45e-07  SA=1.7e-07  SB=5.26e-07  NRD=0.426  NRS=0.684  SCA=15.255  SCB=0.017  SCC=0.002 
R0 M6:DRN M10:SRC 71.8721 
R1 M10:SRC M8:GATE 200.436 
CC80256 M10:SRC M10:GATE 3.589e-17
CC80251 M10:SRC M14:GATE 2.08e-18
CC80226 M10:SRC M9:GATE 9.47e-18
CC80280 M10:SRC M8:DRN 4.398e-17
CC80302 M10:SRC N_9:1 8.41e-18
CC80265 M10:SRC M6:GATE 1.639e-17
CC80332 M10:SRC M8:SRC 3.288e-17
CC80259 M10:SRC A1 7.91e-18
R2 M4:GATE M8:GATE 259.701 
R3 M8:GATE M6:DRN 205.785 
CC80253 M8:GATE M14:GATE 6.25e-18
CC80246 M8:GATE M3:GATE 2.52e-18
CC80356 M8:GATE M4:SRC 1.171e-17
CC80306 M8:GATE N_9:1 4.48e-18
CC80270 M8:GATE M5:GATE 4.12e-18
CC80283 M8:GATE M8:DRN 3.702e-17
CC80328 M8:GATE M8:SRC 5.42e-18
CC80227 M8:GATE M9:GATE 4.07e-18
CC80336 M8:GATE M8:SRC 3.937e-17
CC80292 M8:GATE M5:SRC 2.08e-18
CC80241 M8:GATE A2 1.44e-18
CC80268 M6:DRN M6:GATE 2.463e-17
CC80263 M6:DRN A1 7.228e-17
CC80339 M4:GATE M8:SRC 1.283e-17
CC80349 M4:GATE M4:SRC 1.2e-18
CC80225 M4:GATE M13:SRC 7.23e-18
CC80247 M4:GATE M3:GATE 2.86e-18
CC80315 M4:GATE N_9:2 1.68e-18
CC80272 M4:GATE M5:GATE 3.75e-18
CC80232 M4:GATE M3:SRC 4.761e-17
CC80360 M4:GATE M4:SRC 2.393e-17
CC80242 M4:GATE A2 8.21e-18
C4 M10:SRC 0 5.195e-17
C5 M8:GATE 0 7.451e-17
C6 M6:DRN 0 1.0627e-16
C7 M4:GATE 0 1.849e-17
R8 M11:SRC Z 30.6736 
R9 Z M2:DRN 15.3128 
CC80362 Z M4:SRC 6.186e-17
CC80321 Z M12:GATE 3.94e-18
CC80345 Z M2:GATE 1.57e-18
CC80312 Z N_9:1 1.519e-17
CC80344 Z M1:GATE 6.22e-18
CC80245 Z A2 1.405e-17
CC80325 Z M11:GATE 1.9e-17
R10 M2:DRN M1:SRC 0.001 
CC80343 M2:DRN M1:GATE 3.976e-17
CC80348 M2:DRN M2:GATE 3.977e-17
CC80311 M2:DRN N_9:1 2.932e-17
R11 M11:SRC M12:DRN 0.001 
CC80319 M11:SRC M12:GATE 2.803e-17
CC80324 M11:SRC M11:GATE 2.798e-17
CC80301 M11:SRC N_9:1 8.64e-18
C12 Z 0 1.5121e-16
C13 M2:DRN 0 7.99e-18
C14 M11:SRC 0 8.03e-18
R15 M13:GATE M3:GATE 570.195 
R16 M3:GATE A2 124.103 
CC80310 M3:GATE N_9:1 5.73e-18
CC80248 M3:GATE M3:SRC 4.06e-18
R17 A2 M13:GATE 149.598 
CC80239 A2 M13:SRC 1.137e-17
CC80313 A2 N_9:1 5.73e-18
CC80243 A2 M3:SRC 9.008e-17
CC80363 A2 M4:SRC 4.072e-17
CC80233 M13:GATE M13:SRC 2.08e-17
CC80318 M13:GATE M12:GATE 5.68e-18
CC80300 M13:GATE N_9:1 2.039e-17
CC80236 M13:GATE M3:SRC 5.46e-18
C18 M3:GATE 0 6.378e-17
C19 A2 0 3.887e-17
C20 M13:GATE 0 9.171e-17
R21 M14:GATE M10:GATE 355.1 
R22 M6:GATE M10:GATE 576.865 
R23 M10:GATE A1 193.755 
CC80326 M10:GATE M8:SRC 3.71e-18
CC80333 M10:GATE M8:SRC 1.88e-18
CC80303 M10:GATE N_9:1 6.38e-18
CC80281 M10:GATE M8:DRN 1.99e-18
CC80257 M10:GATE M9:GATE 1.1e-18
R24 A1 M6:GATE 98.7091 
CC80287 A1 M8:DRN 2.118e-17
CC80262 A1 M7:GATE 1.098e-17
CC80260 A1 M9:GATE 5.65e-18
R25 M6:GATE M5:GATE 332.045 
CC80294 M6:GATE M5:SRC 3.26e-18
CC80267 M6:GATE M7:GATE 4.25e-18
CC80269 M6:GATE M3:SRC 1.375e-17
CC80295 M5:GATE M5:SRC 1.422e-17
CC80289 M5:GATE M5:SRC 4.54e-18
CC80286 M5:GATE M8:DRN 3.38e-18
CC80277 M5:GATE N_8:1 1.88e-18
CC80308 M5:GATE N_9:1 5.04e-18
CC80273 M5:GATE M3:SRC 1.478e-17
CC80359 M5:GATE M4:SRC 1.914e-17
CC80299 M14:GATE N_9:1 2.62e-18
CC80330 M14:GATE M8:SRC 2.22e-17
CC80254 M14:GATE M3:SRC 1.55e-18
CC80250 M14:GATE M13:SRC 1.314e-17
CC80255 M14:GATE M13:SRC 1.12e-18
C26 M10:GATE 0 1.521e-16
C27 A1 0 6.587e-17
C28 M6:GATE 0 1.1709e-16
C29 M5:GATE 0 4.315e-17
C30 M14:GATE 0 5.252e-17
R31 M7:GATE M13:SRC 167.799 
R32 M13:SRC M3:SRC 74.2552 
CC80298 M13:SRC N_9:1 6.948e-17
R33 M3:SRC M7:GATE 164.087 
CC80278 M3:SRC N_8:1 4.57e-18
CC80340 M3:SRC M8:SRC 1.276e-17
CC80296 M3:SRC M5:SRC 3.175e-17
CC80361 M3:SRC M4:SRC 4.39e-18
CC80350 M3:SRC M4:SRC 1.42e-18
R34 M7:GATE M9:GATE 137.8 
CC80307 M7:GATE N_9:1 6.221e-17
CC80275 M7:GATE N_8:1 2.47e-18
CC80284 M7:GATE M8:DRN 5.59e-18
CC80293 M7:GATE M5:SRC 3.637e-17
CC80282 M9:GATE M8:DRN 3.757e-17
C35 M13:SRC 0 9.304e-17
C36 M3:SRC 0 5.16e-18
C37 M7:GATE 0 3.809e-17
C38 M9:GATE 0 5.174e-17
R39 N_8:1 M5:SRC 10.6529 
R40 M5:SRC M8:DRN 60.6027 
CC80337 M5:SRC M8:SRC 6.886e-17
CC80335 M8:DRN M8:SRC 1.39e-18
C41 N_8:1 0 1e-19
C42 M5:SRC 0 2.554e-17
C43 M8:DRN 0 2.11e-18
R44 N_9:2 N_9:3 14.1489 
R45 N_9:3 M4:SRC 30.0617 
R46 M8:SRC M4:SRC 99.3746 
R47 N_9:2 M4:SRC 28.887 
R48 M4:SRC N_9:1 79.3008 
R49 M8:SRC N_9:1 77.2655 
R50 M11:GATE N_9:1 148.359 
R51 M1:GATE N_9:1 150.237 
R52 M12:GATE N_9:1 104.675 
R53 N_9:1 M2:GATE 95.7611 
R54 M1:GATE M11:GATE 715.49 
C55 M4:SRC 0 3.734e-17
C56 N_9:1 0 7.087e-17
C57 M2:GATE 0 2.466e-17
C58 N_9:2 0 2.3e-19
C59 M12:GATE 0 6.988e-17
C60 M1:GATE 0 3.232e-17
C61 M11:GATE 0 8.145e-17
C62 M8:SRC 0 3.062e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
