.SUBCKT BUFFD6 I Z
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.75e-06  SB=4.5e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.49e-06  SB=7.1e-07  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7.4e-14  AS=3.9e-14  PD=1.16e-06  PS=5.9e-07  SA=2.01e-06  SB=1.9e-07  NRD=0.531  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.23e-06  SB=9.7e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.75e-06  SB=4.5e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.7e-07  SB=1.23e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.49e-06  SB=7.1e-07  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7.05e-07  SB=1.475e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.23e-06  SB=9.7e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vdd M15:GATE M15:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.45e-07  SB=1.735e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.7e-07  SB=1.23e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M15:SRC M16:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=9.9e-14  PD=7.2e-07  PS=1.42e-06  SA=1.9e-07  SB=2.01e-06  NRD=2.057  NRS=0.554  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.15e-07  SB=1.495e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.55e-07  SB=1.755e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M7:SRC M8:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=7.4e-14  PD=5.9e-07  PS=1.16e-06  SA=1.9e-07  SB=2.01e-06  NRD=4.141  NRS=0.619  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.2e-07  AD=9.9e-14  AS=5.2e-14  PD=1.42e-06  PS=7.2e-07  SA=2.01e-06  SB=1.9e-07  NRD=0.466  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M12:DRN Z 15.5331 
R1 M10:DRN Z 15.5176 
R2 M2:DRN Z 15.4551 
R3 M4:DRN Z 15.5172 
R4 M6:DRN Z 15.662 
R5 Z M14:DRN 15.7312 
CC77970 Z M15:SRC 3.199e-17
CC77973 Z M4:GATE 1.652e-17
CC77978 Z M3:GATE 1.326e-17
CC77979 Z M2:GATE 1.234e-17
CC77982 Z M1:GATE 3.76e-18
CC77966 Z N_14:4 6.997e-17
CC77963 Z M9:GATE 6.1e-18
CC77960 Z M10:GATE 1.993e-17
CC77957 Z M11:GATE 2.627e-17
CC77954 Z M12:GATE 1.95e-17
CC78001 Z M7:SRC 1.1e-18
CC77987 Z M5:GATE 1.477e-17
CC77951 Z M13:GATE 1.599e-17
CC77946 Z M14:GATE 5.1e-18
CC77938 Z N_14:2 5.87e-18
CC77932 Z N_14:1 6.367e-17
R6 M12:DRN M14:DRN 662.299 
R7 M14:DRN M13:SRC 0.001 
CC77995 M14:DRN M7:SRC 1.33e-18
CC77949 M14:DRN M13:GATE 4.538e-17
CC77945 M14:DRN M14:GATE 4.617e-17
CC77925 M14:DRN N_14:1 1.016e-17
R8 M4:DRN M6:DRN 680.221 
R9 M6:DRN M5:SRC 0.001 
CC77985 M6:DRN M5:GATE 5.1e-18
CC77964 M6:DRN N_14:4 4.079e-17
CC77999 M6:DRN M7:SRC 1.81e-18
CC77990 M6:DRN M6:GATE 1.227e-17
CC77935 M6:DRN N_14:2 1.25e-18
CC77929 M6:DRN N_14:1 5.006e-17
R10 M4:DRN M3:SRC 0.001 
CC77975 M4:DRN M4:GATE 5.07e-18
CC77976 M4:DRN M3:GATE 8.16e-18
CC77940 M4:DRN N_14:3 5.818e-17
CC77936 M4:DRN N_14:2 2.06e-17
CC77930 M4:DRN N_14:1 1.592e-17
R11 M2:DRN M1:SRC 0.001 
CC77981 M2:DRN M2:GATE 5.02e-18
CC77983 M2:DRN M1:GATE 1.819e-17
CC77941 M2:DRN N_14:3 2.09e-18
CC77937 M2:DRN N_14:2 6.968e-17
CC77931 M2:DRN N_14:1 1.615e-17
R12 M10:DRN M9:SRC 0.001 
CC77961 M10:DRN M9:GATE 4.625e-17
CC77959 M10:DRN M10:GATE 4.503e-17
CC77927 M10:DRN N_14:1 1.035e-17
R13 M12:DRN M11:SRC 0.001 
CC77955 M12:DRN M11:GATE 4.5e-17
CC77953 M12:DRN M12:GATE 4.52e-17
CC77926 M12:DRN N_14:1 1.01e-17
C14 Z 0 3.2979e-16
C15 M14:DRN 0 1.035e-17
C16 M6:DRN 0 8.66e-18
C17 M4:DRN 0 8.73e-18
C18 M2:DRN 0 8.26e-18
C19 M10:DRN 0 1.07e-17
C20 M12:DRN 0 8.44e-18
R21 I M15:GATE 440.773 
R22 M7:GATE M15:GATE 727.844 
R23 M15:GATE I:1 239.191 
CC77994 M15:GATE M7:SRC 7.56e-18
CC77944 M15:GATE M14:GATE 7.09e-18
CC77969 M15:GATE M15:SRC 4.732e-17
R24 M8:GATE I:1 94.0755 
R25 I I:1 38.8793 
R26 M7:GATE I:1 202.173 
R27 I:1 M16:GATE 111.3 
CC77972 I:1 M15:SRC 2.982e-17
CC77934 I:1 N_14:1 6.12e-18
CC78003 I:1 M7:SRC 4.948e-17
CC77993 M16:GATE M7:SRC 4.56e-18
CC77968 M16:GATE M15:SRC 4.598e-17
R28 M7:GATE I 372.557 
CC77989 M7:GATE M6:GATE 1.55e-18
CC77928 M7:GATE N_14:1 4.67e-18
CC77998 M7:GATE M7:SRC 1.324e-17
CC77992 I M6:GATE 2.81e-18
CC77971 I M15:SRC 7.825e-17
CC78002 I M7:SRC 1.647e-17
CC77997 M8:GATE M7:SRC 4.271e-17
C29 M15:GATE 0 8.327e-17
C30 I:1 0 4.353e-17
C31 M16:GATE 0 7.307e-17
C32 M7:GATE 0 6.126e-17
C33 I 0 6.317e-17
C34 M8:GATE 0 2.258e-17
R35 M14:GATE N_14:1 111.3 
R36 M15:SRC N_14:1 76.7488 
R37 M7:SRC N_14:1 75.9761 
R38 M6:GATE N_14:1 80.8704 
R39 N_14:1 N_14:4 19.1085 
R40 N_14:3 N_14:4 21.2313 
R41 M15:SRC N_14:4 77.8106 
R42 M7:SRC N_14:4 77.0264 
R43 M13:GATE N_14:4 111.3 
R44 N_14:4 M5:GATE 82.3623 
R45 M7:SRC M15:SRC 53.6344 
R46 M2:GATE N_14:2 94.0755 
R47 M10:GATE N_14:2 111.3 
R48 M11:GATE N_14:2 275.689 
R49 M3:GATE N_14:2 233.022 
R50 N_14:3 N_14:2 60.2341 
R51 M9:GATE N_14:2 164.389 
R52 N_14:2 M1:GATE 138.947 
R53 M1:GATE M9:GATE 635.948 
R54 M4:GATE N_14:3 94.0755 
R55 M12:GATE N_14:3 111.3 
R56 M11:GATE N_14:3 275.689 
R57 N_14:3 M3:GATE 233.022 
R58 M3:GATE M11:GATE 1066.52 
C59 M14:GATE 0 7.138e-17
C60 N_14:1 0 1.3228e-16
C61 N_14:4 0 2.257e-17
C62 M5:GATE 0 3.151e-17
C63 M13:GATE 0 4.883e-17
C64 M6:GATE 0 4.283e-17
C65 M7:SRC 0 1.1037e-16
C66 M15:SRC 0 8.69e-18
C67 N_14:2 0 2.268e-17
C68 M1:GATE 0 5.773e-17
C69 M9:GATE 0 9.817e-17
C70 N_14:3 0 8.96e-18
C71 M3:GATE 0 3.835e-17
C72 M11:GATE 0 4.717e-17
C73 M12:GATE 0 4.314e-17
C74 M10:GATE 0 5.019e-17
C75 M2:GATE 0 4.143e-17
C76 M4:GATE 0 2.925e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
