.SUBCKT AOI21D1 A1 A2 B ZN
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4.1e-14  PD=5.9e-07  PS=6e-07  SA=4.3e-07  SB=4.6e-07  NRD=4.183  NRS=2.587  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.97e-07  AD=7.8e-14  AS=3.9e-14  PD=1.18e-06  PS=5.9e-07  SA=6.9e-07  SB=2e-07  NRD=1.346  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M1:SRC M3:GATE vss vss nch L=6e-08 W=3.9e-07  AD=4.1e-14  AS=6.2e-14  PD=6e-07  PS=1.1e-06  SA=1.6e-07  SB=7.3e-07  NRD=2.587  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE M4:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.3e-07  SB=4.6e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 M4:DRN M5:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=1.04e-13  PD=7.2e-07  PS=1.44e-06  SA=6.9e-07  SB=2e-07  NRD=2.099  NRS=1.435  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE M6:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.8e-14  PD=7.2e-07  PS=1.38e-06  SA=1.7e-07  SB=7.2e-07  NRD=2.099  NRS=0.538  SCA=9.643  SCB=0.01  SCC=0.000823 
CC90782 M1:SRC A1 1.05e-18
R0 A1 M4:GATE 142.907 
R1 M4:GATE M1:GATE 544.696 
CC90749 M4:GATE M4:DRN 2.955e-17
CC90750 M4:GATE M4:SRC 2.807e-17
CC90751 M4:GATE ZN 5.07e-18
CC90752 M4:GATE B 1.45e-18
CC90748 M4:GATE M5:GATE 6.69e-18
CC90773 M4:GATE A2 1.722e-17
CC90747 M4:GATE M6:SRC 4.54e-18
CC90767 M4:GATE M6:GATE 7.44e-18
R2 M1:GATE A1 125.114 
CC90762 M1:GATE ZN 4.1e-18
CC90763 M1:GATE B 3.98e-18
CC90780 M1:GATE M3:GATE 4.01e-18
CC90760 M1:GATE M4:SRC 1.74e-18
CC90761 M1:GATE M2:GATE 3.91e-18
CC90775 M1:GATE A2 4.99e-18
CC90753 A1 M5:GATE 6.84e-18
CC90769 A1 M6:GATE 1.62e-18
CC90778 A1 M3:GATE 8.13e-18
CC90759 A1 B 4.512e-17
CC90758 A1 ZN 3.875e-17
CC90757 A1 M2:GATE 1.148e-17
CC90777 A1 A2 2.307e-17
CC90756 A1 M2:SRC 3.029e-17
CC90755 A1 M4:SRC 4.45e-18
CC90754 A1 M4:DRN 2.7e-18
C3 M4:GATE 0 3.383e-17
C4 M1:GATE 0 3.776e-17
C5 A1 0 1.175e-17
R6 ZN M4:SRC 31.4775 
R7 M4:SRC M6:DRN 0.001 
CC90766 M4:SRC M6:GATE 2.832e-17
CC90732 M4:SRC M4:DRN 5.81e-18
R8 M1:DRN M2:SRC 0.001 
R9 M2:SRC ZN 30.8709 
CC90740 M2:SRC M5:GATE 2.34e-18
CC90744 M2:SRC B 3.234e-17
CC90741 ZN M5:GATE 9.08e-18
CC90745 ZN B 7.284e-17
CC90746 ZN M2:GATE 1.538e-17
CC90776 ZN A2 6.45e-18
CC90768 ZN M6:GATE 2.27e-18
CC90734 ZN M4:DRN 7.659e-17
C10 M4:SRC 0 4.49e-18
C11 M2:SRC 0 4.97e-18
C12 ZN 0 1.3272e-16
R13 M6:SRC M4:DRN 60.7495 
CC90770 M6:SRC A2 7.89e-18
CC90764 M6:SRC M6:GATE 3.549e-17
CC90779 M6:SRC M3:GATE 2.6e-18
CC90737 M6:SRC M5:GATE 1.45e-18
CC90771 M4:DRN A2 1.755e-17
CC90742 M4:DRN B 5.77e-18
CC90738 M4:DRN M5:GATE 3.346e-17
C14 M6:SRC 0 9.924e-17
C15 M4:DRN 0 7.17e-18
R16 M2:GATE B 125.114 
R17 B M5:GATE 142.907 
R18 M5:GATE M2:GATE 544.696 
C19 B 0 2.836e-17
C20 M5:GATE 0 7.583e-17
C21 M2:GATE 0 4.705e-17
R22 M3:GATE A2 120.972 
R23 A2 M6:GATE 139.043 
R24 M6:GATE M3:GATE 504.541 
C25 A2 0 6.752e-17
C26 M6:GATE 0 4.757e-17
C27 M3:GATE 0 5.227e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
