.SUBCKT BUFFD1 I Z
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=2.02e-07  AD=3.7e-14  AS=2.3e-14  PD=7.7e-07  PS=3.93e-07  SA=1.9e-07  SB=4.25e-07  NRD=1.02  NRS=0.611  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=6.4e-14  AS=4.5e-14  PD=1.11e-06  PS=7.87e-07  SA=2.32e-07  SB=1.65e-07  NRD=0.474  NRS=8.098  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=4.5e-14  AS=3e-14  PD=8.7e-07  PS=4.8e-07  SA=1.75e-07  SB=4.25e-07  NRD=0.754  NRS=0.469  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM4 M4:DRN M4:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=8.6e-14  AS=6.1e-14  PD=1.37e-06  PS=9.6e-07  SA=2.3e-07  SB=1.65e-07  NRD=0.433  NRS=7.19  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M4:DRN Z 15.4262 
R1 Z M2:DRN 15.2536 
CC77757 Z M1:DRN 3.782e-17
CC77754 Z M2:GATE 1.107e-17
CC77752 Z M3:DRN 7.93e-18
CC77751 Z M4:GATE 2.875e-17
CC77756 M2:DRN M1:DRN 4.356e-17
CC77753 M2:DRN M2:GATE 6.9e-18
CC77755 M4:DRN M1:DRN 1.59e-18
CC77750 M4:DRN M4:GATE 4.763e-17
C2 Z 0 1.1311e-16
C3 M2:DRN 0 2.594e-17
C4 M4:DRN 0 2.719e-17
R5 M1:GATE I 142.332 
R6 I M3:GATE 178.301 
CC77761 I M4:GATE 1.309e-17
CC77762 I M3:DRN 9.334e-17
CC77763 I M2:GATE 5.1e-18
CC77764 I M1:DRN 1.554e-17
R7 M3:GATE M1:GATE 832.919 
CC77758 M3:GATE M4:GATE 6.39e-18
CC77759 M3:GATE M3:DRN 2.928e-17
CC77760 M3:GATE M1:DRN 4.01e-18
CC77767 M1:GATE M1:DRN 3.266e-17
CC77765 M1:GATE M3:DRN 1.51e-18
CC77766 M1:GATE M2:GATE 1.54e-18
C8 I 0 4.632e-17
C9 M3:GATE 0 9.516e-17
C10 M1:GATE 0 5.087e-17
R11 M2:GATE M1:DRN 299.101 
R12 M3:DRN M1:DRN 76.914 
R13 M1:DRN M4:GATE 362.546 
R14 M2:GATE M4:GATE 392.325 
R15 M4:GATE M3:DRN 363.682 
R16 M3:DRN M2:GATE 300.039 
C17 M1:DRN 0 7.563e-17
C18 M4:GATE 0 8.736e-17
C19 M3:DRN 0 7.607e-17
C20 M2:GATE 0 9.511e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
