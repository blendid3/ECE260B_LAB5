.SUBCKT DFCSNQD1 D CP CDN SDN Q
MMM20 M20:DRN M20:GATE vdd vdd pch L=6e-08 W=1.55e-07  AD=2.6e-14  AS=2e-14  PD=6.5e-07  PS=4.15e-07  SA=1.75e-07  SB=6.2e-07  NRD=1.195  NRS=0.955  SCA=14.652  SCB=0.018  SCC=0.001 
MMM21 M21:DRN M21:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=4.1e-14  AS=2.3e-14  PD=8.4e-07  PS=4.4e-07  SA=4e-07  SB=1.58e-07  NRD=0.698  NRS=12.397  SCA=5.267  SCB=0.005  SCC=7.585e-05 
MMM22 M22:DRN M22:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=4.2e-14  AS=2.3e-14  PD=8.4e-07  PS=4.4e-07  SA=1.6e-07  SB=3.98e-07  NRD=0.704  NRS=12.397  SCA=5.267  SCB=0.005  SCC=7.585e-05 
MMM23 M23:DRN M23:GATE M23:SRC vdd pch L=6e-08 W=1.53e-07  AD=2.6e-14  AS=1.7e-14  PD=6.5e-07  PS=3.35e-07  SA=4.25e-07  SB=1.75e-07  NRD=1.195  NRS=0.755  SCA=20.527  SCB=0.023  SCC=0.003 
MMM24 M24:DRN M24:GATE M23:SRC vdd pch L=6e-08 W=2.8e-07  AD=4.4e-14  AS=3.1e-14  PD=8.9e-07  PS=6.25e-07  SA=1.55e-07  SB=2.28e-07  NRD=0.66  NRS=14.264  SCA=14.603  SCB=0.016  SCC=0.002 
MMM25 vdd M25:GATE M25:SRC vdd pch L=6e-08 W=4.82e-07  AD=6.7e-14  AS=4.8e-14  PD=1.36e-06  PS=6.8e-07  SA=4.96e-07  SB=1.34e-07  NRD=0.524  NRS=2.258  SCA=10.228  SCB=0.011  SCC=0.0008915 
MMM26 M25:SRC M26:GATE vdd vdd pch L=6e-08 W=4.84e-07  AD=4.8e-14  AS=6.4e-14  PD=6.8e-07  PS=1.329e-06  SA=2e-07  SB=3.97e-07  NRD=2.258  NRS=0.731  SCA=7.816  SCB=0.008  SCC=0.0004769 
MMM27 M19:DRN M27:GATE vdd vdd pch L=6e-08 W=1.58e-07  AD=2.4e-14  AS=2e-14  PD=5.18e-07  PS=4.15e-07  SA=1.3e-07  SB=2.5e-07  NRD=1.072  NRS=0.955  SCA=3.346  SCB=0.002  SCC=4.515e-06 
MMM28 M19:SRC M28:GATE M28:SRC vdd pch L=6e-08 W=4.95e-07  AD=5.9e-14  AS=3.5e-14  PD=1.019e-06  PS=6.35e-07  SA=3.3e-07  SB=1.91e-07  NRD=10.371  NRS=14.773  SCA=8.408  SCB=0.009  SCC=0.0005868 
MMM29 M28:SRC M29:GATE vdd vdd pch L=6e-08 W=4.99e-07  AD=3.5e-14  AS=6.4e-14  PD=6.35e-07  PS=1.25e-06  SA=1.3e-07  SB=4.12e-07  NRD=14.773  NRS=1.814  SCA=8.408  SCB=0.009  SCC=0.0005868 
MMM10 M10:DRN M10:GATE M10:SRC vss nch L=6e-08 W=1.5e-07  AD=1.3e-14  AS=1.3e-14  PD=3.2e-07  PS=3.2e-07  SA=6.85e-07  SB=1.356e-06  NRD=22.667  NRS=22.667  SCA=20.648  SCB=0.023  SCC=0.003 
MMM11 M11:DRN M11:GATE M11:SRC vss nch L=6e-08 W=3.94e-07  AD=3.8e-14  AS=4.4e-14  PD=6.62e-07  PS=8.52e-07  SA=2.71e-07  SB=2.17e-07  NRD=8.254  NRS=10.891  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=2.1e-07  AD=3.9e-14  AS=1.7e-14  PD=7.9e-07  PS=3.7e-07  SA=1.85e-07  SB=8.95e-07  NRD=0.935  NRS=19.037  SCA=17.402  SCB=0.019  SCC=0.002 
MMM12 M8:SRC M12:GATE M12:SRC vss nch L=6.1e-08 W=2.32e-07  AD=2.5e-14  AS=2.5e-14  PD=4.81e-07  PS=5.21e-07  SA=5.54e-07  SB=2.7e-07  NRD=5.114  NRS=11.621  SCA=16.515  SCB=0.019  SCC=0.002 
MMM2 M2:DRN M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=7e-14  AS=2.9e-14  PD=1.14e-06  PS=5.4e-07  SA=5.61e-07  SB=1.8e-07  NRD=0.508  NRS=11.783  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M11:DRN vss nch L=6e-08 W=3.1e-07  AD=5.3e-14  AS=3e-14  PD=9.6e-07  PS=5.18e-07  SA=1.75e-07  SB=3.78e-07  NRD=0.676  NRS=1.015  SCA=7.268  SCB=0.008  SCC=0.0002566 
MMM3 M1:SRC M3:GATE vss vss nch L=6e-08 W=2.17e-07  AD=1.7e-14  AS=2.8e-14  PD=3.7e-07  PS=4.31e-07  SA=4.05e-07  SB=6.75e-07  NRD=19.037  NRS=0.625  SCA=17.402  SCB=0.019  SCC=0.002 
MMM14 M12:SRC M14:GATE M14:SRC vss nch L=6e-08 W=1.55e-07  AD=1.7e-14  AS=2.6e-14  PD=3.39e-07  PS=6.5e-07  SA=9.56e-07  SB=1.75e-07  NRD=0.746  NRS=1.195  SCA=20.622  SCB=0.023  SCC=0.003 
MMM4 vss M4:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=5.1e-14  AS=2.9e-14  PD=7.99e-07  PS=5.4e-07  SA=3.03e-07  SB=3.9e-07  NRD=3.924  NRS=11.783  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 M10:DRN M15:GATE vss vss nch L=6e-08 W=1.59e-07  AD=1.3e-14  AS=2.1e-14  PD=3.2e-07  PS=3.83e-07  SA=9.2e-07  SB=1.124e-06  NRD=22.667  NRS=1.048  SCA=20.648  SCB=0.023  SCC=0.003 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.2e-14  AS=5.3e-14  PD=1.1e-06  PS=1.05e-06  SA=1.35e-07  SB=1.6e-07  NRD=0.462  NRS=1.581  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M11:SRC M16:GATE M10:SRC vss nch L=6e-08 W=1.56e-07  AD=1.7e-14  AS=1.3e-14  PD=3.28e-07  PS=3.2e-07  SA=4.48e-07  SB=1.588e-06  NRD=0.762  NRS=22.667  SCA=20.648  SCB=0.023  SCC=0.003 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=2.04e-07  AD=3.4e-14  AS=1.8e-14  PD=7.4e-07  PS=3.75e-07  SA=4.15e-07  SB=1.75e-07  NRD=0.947  NRS=14.653  SCA=8.121  SCB=0.009  SCC=0.0003028 
MMM17 vdd M17:GATE M17:SRC vdd pch L=6e-08 W=3.54e-07  AD=4.5e-14  AS=3.5e-14  PD=9.6e-07  PS=5.5e-07  SA=1.35e-07  SB=1.38e-06  NRD=1.551  NRS=3.039  SCA=12.653  SCB=0.014  SCC=0.001 
MMM7 M7:DRN M7:GATE vss vss nch L=6e-08 W=2.04e-07  AD=3.4e-14  AS=1.8e-14  PD=7.4e-07  PS=3.75e-07  SA=1.75e-07  SB=4.15e-07  NRD=0.947  NRS=14.653  SCA=8.121  SCB=0.009  SCC=0.0003028 
MMM18 M17:SRC M18:GATE vdd vdd pch L=6e-08 W=3.55e-07  AD=3.5e-14  AS=4.1e-14  PD=5.5e-07  PS=5.91e-07  SA=3.96e-07  SB=1.12e-06  NRD=3.039  NRS=0.598  SCA=12.653  SCB=0.014  SCC=0.001 
MMM8 M8:DRN M8:GATE M8:SRC vss nch L=6e-08 W=2.12e-07  AD=1.5e-14  AS=2.3e-14  PD=3.5e-07  PS=4.39e-07  SA=8.38e-07  SB=4.34e-07  NRD=24.729  NRS=0.538  SCA=12.705  SCB=0.015  SCC=0.001 
MMM19 M19:DRN M19:GATE M19:SRC vdd pch L=6e-08 W=1.87e-07  AD=2.9e-14  AS=2.1e-14  PD=6.22e-07  PS=3.71e-07  SA=5.9e-07  SB=1.8e-07  NRD=0.9  NRS=0.667  SCA=6.102  SCB=0.006  SCC=0.0001158 
MMM9 M8:DRN M9:GATE vss vss nch L=6e-08 W=2.18e-07  AD=1.5e-14  AS=2.9e-14  PD=3.5e-07  PS=5.37e-07  SA=5.23e-07  SB=6.79e-07  NRD=24.729  NRS=0.881  SCA=14.662  SCB=0.017  SCC=0.001 
MMM30 M30:DRN M30:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=9.5e-14  PD=1.36e-06  PS=8.85e-07  SA=1.134e-06  SB=1.6e-07  NRD=0.427  NRS=0.639  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM31 vdd M31:GATE M31:SRC vdd pch L=6e-08 W=5.22e-07  AD=9.5e-14  AS=5.2e-14  PD=8.85e-07  PS=7.2e-07  SA=6.71e-07  SB=5.85e-07  NRD=0.639  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM32 M31:SRC M32:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.1e-14  PD=7.2e-07  PS=8.79e-07  SA=3.43e-07  SB=8.45e-07  NRD=2.099  NRS=3.178  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M5:DRN Q 15.2649 
CC66602 M5:DRN N_17:1 4.049e-17
CC66641 M5:DRN M5:GATE 1.029e-17
R1 Q M30:DRN 15.4128 
CC66606 Q N_17:1 7.67e-17
CC66613 Q M30:GATE 9.78e-18
CC66644 Q M5:GATE 5.07e-18
CC66651 Q M2:DRN 3.035e-17
CC66596 M30:DRN N_17:1 5.31e-18
CC66612 M30:DRN M30:GATE 4.643e-17
C2 M5:DRN 0 1.677e-17
C3 Q 0 8.007e-17
C4 M30:DRN 0 1.905e-17
CC66427 M1:SRC CDN:1 1.18e-18
CC66670 M10:SRC N_35:1 1.41e-18
CC66586 M11:DRN M13:GATE 3.25e-18
CC66425 M11:DRN D 1.6e-18
R5 M25:GATE M17:GATE 536.624 
R6 M1:GATE M17:GATE 357.824 
R7 M17:GATE SDN 130.423 
CC66408 M17:GATE M23:DRN 1.299e-17
CC66409 M17:GATE M17:SRC 2.065e-17
CC66410 M17:GATE M1:DRN 2.1e-18
CC66633 M17:GATE M3:GATE 1.5e-18
CC66625 M17:GATE M18:GATE 1.79e-18
CC66600 M17:GATE N_17:1 6.17e-18
R8 SDN M1:GATE 99.9317 
CC66478 SDN M23:GATE 2.27e-18
CC66411 SDN M23:DRN 2.07e-18
CC66412 SDN M17:SRC 9.725e-17
CC66414 SDN M1:DRN 1.37e-17
CC66637 SDN M3:GATE 1.51e-17
CC66628 SDN M18:GATE 3.01e-18
CC66415 M1:GATE M23:DRN 3.96e-18
CC66416 M1:GATE M1:DRN 2.329e-17
CC66464 M1:GATE N_24:1 6.19e-18
CC66635 M1:GATE M3:GATE 6.49e-18
R9 M25:GATE M8:GATE 182.85 
CC66678 M25:GATE M24:DRN 3.54e-18
CC66418 M25:GATE M23:DRN 1.55e-18
CC66420 M25:GATE M11:SRC 4.13e-18
CC66485 M25:GATE M12:GATE 3.94e-18
CC66417 M25:GATE M26:GATE 8.12e-18
CC66721 M25:GATE M8:SRC 9.46e-18
CC66657 M25:GATE N_35:1 5.14e-18
CC66470 M25:GATE M23:GATE 1.25e-18
CC66597 M25:GATE N_17:1 5.12e-18
CC66706 M25:GATE M25:SRC 3.146e-17
CC66684 M8:GATE M24:DRN 2.04e-18
CC66424 M8:GATE M9:GATE 2.622e-17
CC66463 M8:GATE N_24:1 9.09e-18
CC66672 M8:GATE N_35:1 7.68e-18
CC66727 M8:GATE M8:SRC 2.212e-17
C10 M17:GATE 0 9.61e-17
C11 SDN 0 2.123e-17
C12 M1:GATE 0 1.663e-17
C13 M25:GATE 0 2.2975e-16
C14 M8:GATE 0 1.385e-17
R15 M1:DRN M17:SRC 125.577 
R16 M14:SRC M17:SRC 125.085 
R17 M17:SRC M23:DRN 118.617 
CC66431 M17:SRC N_28:1 1.782e-17
CC66599 M17:SRC N_17:1 2.15e-17
CC66624 M17:SRC M18:GATE 1.348e-17
R18 M1:DRN M23:DRN 122.983 
R19 M23:DRN M14:SRC 122.501 
CC66391 M23:DRN CDN 1.13e-17
CC66393 M23:DRN CDN:1 3.7e-18
CC66472 M23:DRN M23:GATE 3.474e-17
CC66430 M23:DRN N_28:1 4.478e-17
CC66486 M23:DRN M12:GATE 1.11e-18
CC66623 M23:DRN M18:GATE 1.22e-18
CC66439 M23:DRN M23:SRC 1.49e-18
CC66454 M23:DRN N_24:1 1.172e-17
CC66531 M23:DRN M14:GATE 2.73e-18
R20 M14:SRC M1:DRN 117.925 
CC66432 M14:SRC N_28:1 4.964e-17
CC66488 M14:SRC M12:GATE 1.71e-18
CC66397 M14:SRC CDN:1 1.96e-18
CC66458 M14:SRC N_24:1 7.436e-17
CC66440 M14:SRC M23:SRC 1.14e-18
CC66532 M14:SRC M14:GATE 2.196e-17
CC66475 M14:SRC M23:GATE 5.34e-18
CC66527 M14:SRC M24:GATE 1.001e-17
CC66491 M1:DRN M12:GATE 2.48e-18
CC66465 M1:DRN N_24:1 1.377e-17
CC66605 M1:DRN N_17:1 3.56e-18
CC66434 M1:DRN N_28:1 6.299e-17
CC66400 M1:DRN CDN:1 5.37e-18
C21 M17:SRC 0 9.5e-19
C22 M23:DRN 0 2.113e-17
C23 M14:SRC 0 4.56e-18
C24 M1:DRN 0 3.716e-17
R25 CP M7:GATE 125.306 
R26 M7:GATE M22:GATE 639.968 
CC66571 M7:GATE M22:DRN 1e-18
CC66578 M7:GATE M6:GATE 8.93e-18
CC66517 M7:GATE N_26:1 6.12e-18
CC66593 M7:GATE M7:DRN 2.325e-17
R27 M22:GATE CP 162.973 
CC66544 M22:GATE N_26:1 8.49e-18
CC66568 M22:GATE M22:DRN 2.943e-17
CC66553 M22:GATE M21:GATE 9.75e-18
CC66510 M22:GATE N_26:1 1.192e-17
CC66570 CP M22:DRN 4.53e-18
CC66549 CP N_26:1 2.397e-17
CC66581 CP M6:GATE 4.99e-18
CC66592 CP M7:DRN 1.481e-17
CC66520 CP N_26:1 8.608e-17
C28 M7:GATE 0 2.803e-17
C29 M22:GATE 0 4.187e-17
C30 CP 0 1.927e-17
R31 M9:GATE M19:SRC 240.775 
R32 M11:SRC M19:SRC 76.4371 
R33 M19:SRC M26:GATE 432.97 
CC66654 M19:SRC N_35:1 6.182e-17
CC66383 M19:SRC M28:GATE 2.79e-17
CC66541 M19:SRC N_26:1 1.74e-18
CC66560 M19:SRC M19:GATE 1.468e-17
CC66388 M19:SRC M11:GATE 1.94e-18
CC66386 M19:SRC D 4.08e-18
CC66505 M19:SRC N_26:1 5.842e-17
CC66450 M19:SRC N_24:1 9.672e-17
R34 M9:GATE M26:GATE 319.562 
R35 M26:GATE M11:SRC 417.899 
CC66656 M26:GATE N_35:1 7.75e-18
CC66543 M26:GATE N_26:1 4.38e-18
CC66401 M26:GATE M20:GATE 7.01e-18
CC66507 M26:GATE N_26:1 2.85e-18
CC66705 M26:GATE M25:SRC 2.105e-17
CC66695 M26:GATE M27:GATE 1.1e-18
CC66451 M26:GATE N_24:1 3.844e-17
R36 M11:SRC M9:GATE 232.391 
CC66664 M11:SRC N_35:1 8.05e-18
CC66515 M11:SRC N_26:1 1.58e-18
CC66382 M11:SRC M19:DRN 1.912e-17
CC66381 M11:SRC M20:DRN 1.965e-17
CC66564 M11:SRC M19:GATE 7.26e-18
CC66406 M11:SRC M15:GATE 1.731e-17
CC66404 M11:SRC M20:GATE 5.73e-18
CC66494 M11:SRC M16:GATE 3.885e-17
CC66389 M11:SRC M11:GATE 4.46e-18
CC66497 M11:SRC M16:GATE 1.64e-18
CC66387 M11:SRC D 9.495e-17
CC66385 M11:SRC M28:GATE 5.04e-18
CC66708 M11:SRC M25:SRC 1.404e-17
CC66456 M11:SRC N_24:1 8.43e-18
CC66460 M11:SRC N_24:1 5.06e-18
CC66722 M11:SRC M8:SRC 1e-18
CC66716 M11:SRC M10:GATE 6.2e-18
CC66671 M9:GATE N_35:1 5.771e-17
CC66398 M9:GATE CDN:1 1.07e-18
CC66718 M9:GATE M10:GATE 2.84e-18
CC66462 M9:GATE N_24:1 1.85e-18
C37 M19:SRC 0 8.1e-18
C38 M26:GATE 0 4.273e-17
C39 M11:SRC 0 1.25e-17
C40 M9:GATE 0 2.473e-17
R41 M20:DRN M19:DRN 60.6736 
CC66402 M20:DRN M20:GATE 3.179e-17
CC66405 M20:DRN M15:GATE 1.37e-18
CC66512 M20:DRN N_26:1 5.57e-18
CC66698 M20:DRN M27:GATE 3.413e-17
CC66661 M20:DRN N_35:1 5.751e-17
CC66506 M19:DRN N_26:1 2.55e-18
CC66513 M19:DRN N_26:1 6.33e-17
CC66403 M19:DRN M20:GATE 3.56e-18
CC66563 M19:DRN M19:GATE 3.442e-17
CC66546 M19:DRN N_26:1 3.43e-18
CC66714 M19:DRN M10:GATE 4.51e-18
CC66662 M19:DRN N_35:1 1.32e-18
CC66700 M19:DRN M27:GATE 2.306e-17
C42 M20:DRN 0 1.206e-17
C43 M19:DRN 0 1.53e-17
R44 D M28:GATE 142.349 
R45 M28:GATE M11:GATE 531.699 
CC66480 M28:GATE M29:GATE 2.115e-17
CC66504 M28:GATE N_26:1 5.25e-18
CC66540 M28:GATE N_26:1 3.08e-18
CC66559 M28:GATE M19:GATE 3.79e-18
R46 M11:GATE D 124.105 
CC66498 M11:GATE M16:GATE 2.12e-18
CC66576 M11:GATE M6:GATE 4.27e-18
CC66461 M11:GATE N_24:1 2.383e-17
CC66519 D N_26:1 1.848e-17
CC66467 D N_24:1 6.319e-17
CC66500 D M16:GATE 3.32e-18
CC66589 D M13:GATE 1.261e-17
CC66482 D M29:GATE 8.25e-18
C47 M28:GATE 0 4.265e-17
C48 M11:GATE 0 2.642e-17
C49 D 0 1.228e-17
R50 M15:GATE CDN:1 109.975 
R51 CDN:1 M4:GATE 681.051 
CC66448 CDN:1 M12:SRC 2.33e-18
CC66445 CDN:1 M2:GATE 5.81e-18
CC66730 CDN:1 M8:SRC 2.78e-18
CC66468 CDN:1 N_24:1 3.054e-17
CC66608 CDN:1 N_17:1 1.58e-18
CC66639 CDN:1 M3:GATE 1.09e-18
R52 CDN M4:GATE 120.869 
R53 M4:GATE M32:GATE 534.776 
CC66443 M4:GATE M2:GATE 4.41e-18
CC66603 M4:GATE N_17:1 2.74e-18
CC66634 M4:GATE M3:GATE 1.315e-17
CC66433 M4:GATE N_28:1 1.264e-17
R54 M32:GATE CDN 146.713 
CC66429 M32:GATE N_28:1 1.049e-17
CC66594 M32:GATE N_17:1 3.85e-18
CC66616 M32:GATE M31:SRC 9.71e-18
CC66622 M32:GATE M18:GATE 1.15e-18
CC66438 CDN M31:GATE 1.496e-17
CC66444 CDN M2:GATE 7.32e-18
CC66607 CDN N_17:1 7.54e-18
CC66620 CDN M31:SRC 1.976e-17
CC66629 CDN M18:GATE 9.36e-18
CC66638 CDN M3:GATE 5.13e-18
CC66435 CDN N_28:1 4.052e-17
R55 M20:GATE M15:GATE 129.849 
CC66697 M20:GATE M27:GATE 2.27e-18
CC66660 M20:GATE N_35:1 1.875e-17
CC66665 M15:GATE N_35:1 7.84e-18
CC66457 M15:GATE N_24:1 9.09e-18
CC66717 M15:GATE M10:GATE 5.59e-18
C56 CDN:1 0 3.3898e-16
C57 M4:GATE 0 6.351e-17
C58 M32:GATE 0 4.475e-17
C59 CDN 0 6.478e-17
C60 M20:GATE 0 2.356e-17
C61 M15:GATE 0 4.335e-17
R62 M12:SRC N_28:1 30.9024 
CC66489 M12:SRC M12:GATE 3.553e-17
CC66668 M12:SRC N_35:1 1.85e-18
CC66459 M12:SRC N_24:1 1.24e-18
CC66682 M12:SRC M24:DRN 1.19e-18
CC66533 M12:SRC M14:GATE 3.449e-17
R63 M31:GATE N_28:1 150.789 
R64 M2:GATE N_28:1 123.873 
R65 N_28:1 M23:SRC 29.9999 
CC66731 N_28:1 M8:SRC 1.01e-18
CC66537 N_28:1 M14:GATE 7.64e-18
CC66567 N_28:1 M19:GATE 7.45e-18
CC66469 N_28:1 N_24:1 2.388e-17
CC66609 N_28:1 N_17:1 1.4657e-16
CC66615 N_28:1 M30:GATE 1.79e-18
CC66621 N_28:1 M31:SRC 1.313e-17
CC66630 N_28:1 M18:GATE 6.45e-18
CC66646 N_28:1 M5:GATE 7.55e-18
CC66653 N_28:1 M2:DRN 3.043e-17
CC66720 N_28:1 M10:GATE 4.75e-18
CC66677 N_28:1 N_35:1 5.834e-17
CC66688 N_28:1 M24:DRN 2.93e-18
CC66492 N_28:1 M12:GATE 5.07e-18
CC66522 N_28:1 N_26:1 1.954e-17
CC66529 N_28:1 M24:GATE 3.15e-18
CC66479 N_28:1 M23:GATE 8.5e-18
CC66471 M23:SRC M23:GATE 3.306e-17
CC66508 M23:SRC N_26:1 1.27e-17
CC66523 M23:SRC M24:GATE 2.09e-17
R66 M2:GATE M31:GATE 488.187 
CC66604 M2:GATE N_17:1 5.77e-18
CC66650 M2:GATE M2:DRN 2.691e-17
CC66611 M31:GATE M30:GATE 4.92e-18
CC66617 M31:GATE M31:SRC 2.958e-17
CC66647 M31:GATE M2:DRN 1.82e-18
CC66595 M31:GATE N_17:1 1.943e-17
C67 M12:SRC 0 4.41e-18
C68 N_28:1 0 7.381e-17
C69 M23:SRC 0 9.86e-18
C70 M2:GATE 0 2.121e-17
C71 M31:GATE 0 2.913e-17
R72 M21:DRN N_24:1 30.6279 
R73 M29:GATE N_24:1 178.025 
R74 M6:DRN N_24:1 30.2136 
R75 M23:GATE N_24:1 262.306 
R76 M12:GATE N_24:1 77.9282 
R77 N_24:1 M16:GATE 87.6242 
CC66591 N_24:1 M13:GATE 5.45e-18
CC66675 N_24:1 N_35:1 3.616e-17
CC66719 N_24:1 M10:GATE 5.17e-18
CC66729 N_24:1 M8:SRC 1.031e-17
CC66557 N_24:1 M21:GATE 9.38e-18
CC66536 N_24:1 M14:GATE 5.89e-18
CC66521 N_24:1 N_26:1 1.2076e-16
CC66550 N_24:1 N_26:1 2.28e-18
CC66582 N_24:1 M6:GATE 1.665e-17
R78 M16:GATE M12:GATE 4532.81 
CC66715 M16:GATE M10:GATE 8.03e-18
CC66663 M16:GATE N_35:1 8.18e-18
R79 M12:GATE M23:GATE 3764.08 
CC66683 M12:GATE M24:DRN 2.08e-18
CC66725 M12:GATE M8:SRC 2.078e-17
CC66534 M12:GATE M14:GATE 3.19e-18
CC66669 M12:GATE N_35:1 5.83e-18
CC66528 M12:GATE M24:GATE 2.53e-18
CC66524 M23:GATE M24:GATE 2.01e-18
CC66530 M23:GATE M14:GATE 5.96e-18
CC66518 M6:DRN N_26:1 1.58e-18
CC66579 M6:DRN M6:GATE 3.662e-17
CC66588 M6:DRN M13:GATE 3.1e-18
CC66539 M29:GATE N_26:1 4.44e-18
CC66503 M29:GATE N_26:1 8.24e-18
CC66551 M29:GATE M21:GATE 1.01e-18
CC66572 M29:GATE M6:GATE 3.11e-18
CC66511 M21:DRN N_26:1 1.445e-17
CC66554 M21:DRN M21:GATE 2.076e-17
C80 N_24:1 0 3.2856e-16
C81 M16:GATE 0 2.583e-17
C82 M12:GATE 0 3.065e-17
C83 M23:GATE 0 1.643e-17
C84 M6:DRN 0 1.664e-17
C85 M29:GATE 0 2.384e-17
C86 M21:DRN 0 1.816e-17
R87 M22:DRN N_26:1 30.1961 
R88 M21:GATE N_26:1 165.97 
R89 M7:DRN N_26:1 31.9685 
R90 M6:GATE N_26:1 131.252 
R91 M19:GATE N_26:1 74.6319 
R92 N_26:1 M24:GATE 83.8599 
CC66711 N_26:1 M25:SRC 8.29e-18
CC66710 N_26:1 M25:SRC 1.42e-18
CC66685 N_26:1 M24:DRN 2.913e-17
CC66702 N_26:1 M27:GATE 5.5e-18
CC66703 N_26:1 M27:GATE 6.9e-18
CC66674 N_26:1 N_35:1 9.211e-17
R93 M19:GATE M24:GATE 4599.43 
R94 M24:GATE M14:GATE 134.941 
CC66658 M24:GATE N_35:1 1.29e-18
CC66679 M24:GATE M24:DRN 1.305e-17
CC66667 M14:GATE N_35:1 1.06e-18
CC66699 M19:GATE M27:GATE 2.48e-18
R95 M13:GATE M6:GATE 248.041 
R96 M21:GATE M6:GATE 640.448 
R97 M6:GATE M7:DRN 5293.67 
C98 N_26:1 0 3.8824e-16
C99 M24:GATE 0 3.402e-17
C100 M14:GATE 0 7.04e-18
C101 M19:GATE 0 1.212e-17
C102 M6:GATE 0 8.103e-17
C103 M7:DRN 0 2.116e-17
C104 M21:GATE 0 1.339e-17
C105 M13:GATE 0 8.267e-17
C106 M22:DRN 0 1.465e-17
R107 M30:GATE M5:GATE 499.441 
R108 M2:DRN M5:GATE 1560.25 
R109 M5:GATE N_17:1 131.086 
R110 M31:SRC N_17:1 29.9999 
R111 M30:GATE N_17:1 159.791 
R112 M2:DRN N_17:1 17.3353 
R113 N_17:1 M18:GATE 98.6657 
R114 M18:GATE M3:GATE 148.93 
R115 M2:DRN M30:GATE 1901.91 
C116 M5:GATE 0 3.85e-17
C117 N_17:1 0 2.1579e-16
C118 M18:GATE 0 3.028e-17
C119 M3:GATE 0 3.122e-17
C120 M2:DRN 0 1.157e-17
C121 M30:GATE 0 4.523e-17
C122 M31:SRC 0 6.08e-18
R123 M24:DRN N_35:1 30.3335 
R124 M8:SRC N_35:1 30.4926 
R125 M25:SRC N_35:1 30.5038 
R126 M27:GATE N_35:1 230.835 
R127 N_35:1 M10:GATE 86.6249 
R128 M10:GATE M27:GATE 528.598 
C129 M24:DRN 0 1.65e-17
C130 N_35:1 0 2.255e-17
C131 M10:GATE 0 4.93e-18
C132 M27:GATE 0 3.795e-17
C133 M25:SRC 0 1.033e-17
C134 M8:SRC 0 6.73e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
