.SUBCKT AOI21D0 A1 A2 B ZN
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=2.02e-07  AD=3.9e-14  AS=2e-14  PD=7.9e-07  PS=3.95e-07  SA=7.05e-07  SB=2e-07  NRD=1.534  NRS=8.262  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM2 M1:SRC M2:GATE M2:SRC vss nch L=6e-08 W=1.95e-07  AD=2e-14  AS=2e-14  PD=3.95e-07  PS=4.05e-07  SA=4.45e-07  SB=4.6e-07  NRD=8.262  NRS=5.175  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM3 M2:SRC M3:GATE vss vss nch L=6e-08 W=1.95e-07  AD=2e-14  AS=3.4e-14  PD=4.05e-07  PS=7.4e-07  SA=1.75e-07  SB=7.3e-07  NRD=5.175  NRS=0.947  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM4 vdd M4:GATE M4:SRC vdd pch L=6e-08 W=2.65e-07  AD=5.2e-14  AS=2.6e-14  PD=9.2e-07  PS=4.6e-07  SA=6.9e-07  SB=2e-07  NRD=0.84  NRS=4.054  SCA=4.783  SCB=0.004  SCC=4.893e-05 
MMM5 M4:SRC M5:GATE M5:SRC vdd pch L=6e-08 W=2.6e-07  AD=2.6e-14  AS=2.7e-14  PD=4.6e-07  PS=4.7e-07  SA=4.3e-07  SB=4.6e-07  NRD=4.054  NRS=0.438  SCA=4.783  SCB=0.004  SCC=4.893e-05 
MMM6 M6:DRN M6:GATE M6:SRC vdd pch L=6e-08 W=2.6e-07  AD=2.7e-14  AS=4.2e-14  PD=4.7e-07  PS=8.4e-07  SA=1.6e-07  SB=7.3e-07  NRD=0.438  NRS=0.704  SCA=4.783  SCB=0.004  SCC=4.893e-05 
R0 M4:GATE B 162.469 
R1 B M1:GATE 152.163 
CC90690 B M4:SRC 1.536e-17
CC90708 B A1 6.87e-17
CC90701 B M5:GATE 3.01e-18
CC90713 B M2:GATE 2.76e-18
CC90692 B ZN 5.741e-17
CC90691 B M1:SRC 1.148e-17
R2 M1:GATE M4:GATE 809.079 
CC90706 M1:GATE A1 8.31e-18
CC90695 M1:GATE ZN 4.88e-18
CC90694 M1:GATE M1:SRC 2.197e-17
CC90711 M1:GATE M2:GATE 2.19e-18
CC90689 M4:GATE ZN 1.119e-17
CC90687 M4:GATE M4:SRC 3.012e-17
CC90685 M4:GATE M6:SRC 4.8e-18
CC90704 M4:GATE A1 1.26e-18
CC90696 M4:GATE M5:GATE 3.28e-18
C3 B 0 3.238e-17
C4 M1:GATE 0 4.475e-17
C5 M4:GATE 0 6.657e-17
R6 A1 M2:GATE 152.163 
R7 M2:GATE M5:GATE 809.079 
CC90712 M2:GATE ZN 2.27e-18
CC90710 M2:GATE M1:SRC 2.26e-17
CC90727 M2:GATE M3:GATE 7.44e-18
CC90722 M2:GATE A2 8.6e-18
R8 M5:GATE A1 162.469 
CC90714 M5:GATE M6:GATE 1.067e-17
CC90699 M5:GATE M4:SRC 3.665e-17
CC90700 M5:GATE ZN 1.161e-17
CC90697 M5:GATE M5:SRC 2.999e-17
CC90730 A1 M3:GATE 1.52e-18
CC90725 A1 A2 1.344e-17
CC90719 A1 M6:GATE 1.45e-18
CC90702 A1 M5:SRC 2.8e-18
CC90705 A1 M1:SRC 1.014e-17
CC90703 A1 M4:SRC 7.21e-18
CC90707 A1 ZN 7.28e-17
C9 M2:GATE 0 1.912e-17
C10 M5:GATE 0 2.737e-17
C11 A1 0 1.46e-17
R12 M1:SRC M5:SRC 1156.3 
R13 ZN M5:SRC 33.4366 
R14 M5:SRC M6:DRN 0.001 
CC90715 M5:SRC M6:GATE 2.63e-17
CC90681 M5:SRC M4:SRC 4.39e-18
R15 ZN M1:SRC 31.8247 
CC90718 ZN M6:GATE 7.1e-18
CC90729 ZN M3:GATE 6.44e-18
CC90724 ZN A2 6.737e-17
CC90682 ZN M6:SRC 5.65e-18
CC90683 ZN M4:SRC 5.234e-17
C16 M5:SRC 0 2.185e-17
C17 ZN 0 1.3729e-16
C18 M1:SRC 0 1.631e-17
R19 A2 M6:GATE 158.744 
R20 M6:GATE M3:GATE 763.281 
CC90717 M6:GATE M4:SRC 8.4e-18
CC90716 M6:GATE M6:SRC 2.952e-17
R21 M3:GATE A2 148.34 
CC90726 M3:GATE M6:SRC 1.8e-18
CC90721 A2 M4:SRC 1.416e-17
CC90720 A2 M6:SRC 4.49e-18
C22 M6:GATE 0 3.409e-17
C23 M3:GATE 0 5.225e-17
C24 A2 0 5.871e-17
R25 M6:SRC M4:SRC 61.2938 
C26 M6:SRC 0 1.2531e-16
C27 M4:SRC 0 1.358e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
