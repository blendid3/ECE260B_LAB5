.SUBCKT ND2D0 A1 A2 ZN
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=1.95e-07  AD=3.6e-14  AS=2e-14  PD=7.6e-07  PS=3.95e-07  SA=4.45e-07  SB=1.85e-07  NRD=0.996  NRS=8.24  SCA=5.381  SCB=0.005  SCC=5.849e-05 
MMM2 vss M2:GATE M1:SRC vss nch L=6e-08 W=1.95e-07  AD=3.6e-14  AS=2e-14  PD=7.6e-07  PS=3.95e-07  SA=1.85e-07  SB=4.45e-07  NRD=0.996  NRS=8.24  SCA=5.381  SCB=0.005  SCC=5.849e-05 
MMM3 vdd M3:GATE M3:SRC vdd pch L=6e-08 W=2.6e-07  AD=4.4e-14  AS=2.6e-14  PD=8.6e-07  PS=4.6e-07  SA=4.3e-07  SB=1.7e-07  NRD=0.737  NRS=4.054  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM4 vdd M4:GATE M4:SRC vdd pch L=6e-08 W=2.6e-07  AD=4.4e-14  AS=2.6e-14  PD=8.6e-07  PS=4.6e-07  SA=1.7e-07  SB=4.3e-07  NRD=0.737  NRS=4.054  SCA=4.031  SCB=0.003  SCC=2.015e-05 
R0 M1:GATE A1 144.414 
R1 A1 M3:GATE 187.24 
CC44922 A1 M4:GATE 4.19e-18
CC44928 A1 A2 3.71e-17
CC44932 A1 M2:GATE 3.71e-18
CC44915 A1 M1:DRN 7.78e-18
CC44916 A1 ZN 8.669e-17
CC44914 A1 M3:SRC 1.42e-18
R2 M3:GATE M1:GATE 897.44 
CC44924 M3:GATE A2 1.18e-18
CC44913 M3:GATE ZN 1.146e-17
CC44912 M3:GATE M3:SRC 3.042e-17
CC44920 M3:GATE M4:GATE 2.04e-18
CC44925 M1:GATE A2 1.193e-17
CC44929 M1:GATE M2:GATE 6.09e-18
CC44917 M1:GATE ZN 5.13e-18
CC44918 M1:GATE M1:DRN 2.557e-17
C3 A1 0 3.546e-17
C4 M3:GATE 0 8.776e-17
C5 M1:GATE 0 1.681e-17
R6 M4:SRC M3:SRC 0.001 
R7 M3:SRC ZN 31.2282 
CC44919 M3:SRC M4:GATE 2.97e-17
R8 ZN M1:DRN 30.5301 
CC44927 ZN A2 1.83e-17
CC44921 ZN M4:GATE 7.98e-18
C9 M3:SRC 0 1.551e-17
C10 ZN 0 1.7099e-16
C11 M1:DRN 0 2.171e-17
R12 A2 M4:GATE 181.152 
R13 M4:GATE M2:GATE 871.021 
R14 M2:GATE A2 145.445 
C15 M4:GATE 0 8.317e-17
C16 M2:GATE 0 5.746e-17
C17 A2 0 8.652e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
