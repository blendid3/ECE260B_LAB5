.SUBCKT OR2XD1 A1 A2 Z
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.8e-14  AS=4.9e-14  PD=1.13e-06  PS=6.4e-07  SA=7.8e-07  SB=1.75e-07  NRD=0.496  NRS=0.654  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.97e-07  AD=4.9e-14  AS=4.1e-14  PD=6.4e-07  PS=6e-07  SA=4.7e-07  SB=4.85e-07  NRD=0.654  NRS=2.647  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M2:SRC M3:GATE vss vss nch L=6e-08 W=3.97e-07  AD=4.1e-14  AS=7.8e-14  PD=6e-07  PS=1.18e-06  SA=2e-07  SB=7.55e-07  NRD=2.647  NRS=1.346  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vdd vdd pch L=6e-08 W=5.23e-07  AD=9.1e-14  AS=7.3e-14  PD=1.39e-06  PS=8e-07  SA=7.75e-07  SB=1.75e-07  NRD=0.446  NRS=0.644  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=5.24e-07  AD=7.3e-14  AS=5.2e-14  PD=8e-07  PS=7.2e-07  SA=4.35e-07  SB=5.15e-07  NRD=0.644  NRS=2.009  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M5:SRC M6:GATE M6:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=9.1e-14  PD=7.2e-07  PS=1.39e-06  SA=1.75e-07  SB=7.75e-07  NRD=2.009  NRS=0.446  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M4:DRN Z 15.4724 
CC73648 M4:DRN M6:SRC 1.65e-18
CC73646 M4:DRN M4:GATE 4.785e-17
R1 Z M1:DRN 15.266 
CC73647 Z M4:GATE 5.52e-18
CC73650 Z M6:SRC 8.226e-17
CC73652 Z M1:GATE 1.042e-17
CC73649 M1:DRN M6:SRC 4.097e-17
CC73651 M1:DRN M1:GATE 9.55e-18
C2 M4:DRN 0 3.155e-17
C3 Z 0 1.0225e-16
C4 M1:DRN 0 2.26e-17
R5 M6:SRC M4:GATE 258.825 
R6 M2:SRC M4:GATE 488.309 
R7 M4:GATE M1:GATE 411.537 
CC73657 M4:GATE A2 1.104e-17
CC73655 M4:GATE M5:GATE 4.32e-18
R8 M6:SRC M1:GATE 212.732 
R9 M1:GATE M2:SRC 401.352 
CC73661 M1:GATE M2:GATE 2.65e-18
CC73670 M1:GATE A1 1.501e-17
CC73659 M1:GATE A2 2.13e-18
R10 M2:SRC M6:SRC 54.8362 
CC73658 M2:SRC A2 1.3301e-16
CC73668 M2:SRC A1 4.464e-17
CC73662 M6:SRC M6:GATE 5.591e-17
CC73660 M6:SRC M2:GATE 7.97e-18
CC73672 M6:SRC M3:GATE 6.38e-18
CC73666 M6:SRC A1 2.12e-17
CC73654 M6:SRC M5:GATE 1.711e-17
C11 M4:GATE 0 8.975e-17
C12 M1:GATE 0 7.33e-17
C13 M2:SRC 0 3.222e-17
C14 M6:SRC 0 1.21e-16
R15 A2 M5:GATE 145.493 
R16 M5:GATE M2:GATE 525.751 
CC73667 M5:GATE A1 1.098e-17
CC73663 M5:GATE M6:GATE 1.374e-17
R17 M2:GATE A2 119.582 
CC73669 M2:GATE A1 1.57e-18
CC73673 M2:GATE M3:GATE 6.33e-18
CC73665 A2 M6:GATE 4.12e-18
CC73674 A2 M3:GATE 3.71e-18
CC73671 A2 A1 2.911e-17
C18 M5:GATE 0 7.57e-17
C19 M2:GATE 0 5.296e-17
C20 A2 0 2.469e-17
R21 M3:GATE M6:GATE 511.383 
R22 M6:GATE A1 144.734 
R23 A1 M3:GATE 118.637 
C24 M6:GATE 0 5.412e-17
C25 A1 0 6.281e-17
C26 M3:GATE 0 4.546e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
