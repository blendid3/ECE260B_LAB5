.SUBCKT BUFFD0 I Z
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=1.95e-07  AD=3.5e-14  AS=2e-14  PD=7.5e-07  PS=3.95e-07  SA=1.8e-07  SB=4.35e-07  NRD=0.972  NRS=8.262  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=1.95e-07  AD=3.4e-14  AS=2e-14  PD=7.4e-07  PS=3.95e-07  SA=4.4e-07  SB=1.75e-07  NRD=0.947  NRS=8.262  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM3 M3:DRN M3:GATE vdd vdd pch L=6e-08 W=2.6e-07  AD=4.5e-14  AS=2.6e-14  PD=8.7e-07  PS=4.6e-07  SA=1.75e-07  SB=4.25e-07  NRD=0.754  NRS=4.054  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM4 M4:DRN M4:GATE vdd vdd pch L=6e-08 W=2.6e-07  AD=4.3e-14  AS=2.6e-14  PD=8.5e-07  PS=4.6e-07  SA=4.35e-07  SB=1.65e-07  NRD=0.72  NRS=4.054  SCA=4.031  SCB=0.003  SCC=2.015e-05 
R0 M2:DRN Z 30.411 
CC77739 M2:DRN M1:DRN 9.41e-18
CC77736 M2:DRN M2:GATE 2.254e-17
R1 Z M4:DRN 30.5787 
CC77740 Z M1:DRN 7.867e-17
CC77735 Z M4:GATE 1.194e-17
CC77737 Z M2:GATE 4.91e-18
CC77734 M4:DRN M4:GATE 2.975e-17
C2 M2:DRN 0 2.282e-17
C3 Z 0 1.1223e-16
C4 M4:DRN 0 2.423e-17
R5 M1:GATE M3:GATE 825.382 
R6 M3:GATE I 186.295 
CC77741 M3:GATE M4:GATE 1.277e-17
CC77742 M3:GATE M3:DRN 2.957e-17
CC77743 M3:GATE M1:DRN 5.47e-18
R7 I M1:GATE 135.469 
CC77744 I M3:DRN 8.383e-17
CC77745 I M2:GATE 2.505e-17
CC77746 I M1:DRN 1.964e-17
CC77747 M1:GATE M2:GATE 1.44e-18
CC77748 M1:GATE M3:DRN 1.3e-18
CC77749 M1:GATE M1:DRN 3.164e-17
C8 M3:GATE 0 8.082e-17
C9 I 0 3.792e-17
C10 M1:GATE 0 5.033e-17
R11 M4:GATE M1:DRN 433.698 
R12 M3:DRN M1:DRN 74.2159 
R13 M1:DRN M2:GATE 348.937 
R14 M4:GATE M2:GATE 617.907 
R15 M2:GATE M3:DRN 349.887 
R16 M3:DRN M4:GATE 434.884 
C17 M1:DRN 0 6.987e-17
C18 M2:GATE 0 6.223e-17
C19 M3:DRN 0 9.528e-17
C20 M4:GATE 0 9.486e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
