.SUBCKT INVD20 I ZN
MMM20 vss M20:GATE M20:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.6e-07  SB=5.04e-06  NRD=0.567  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM21 vdd M21:GATE M21:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=5.04e-06  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=4.78e-06  SB=4.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 vdd M23:GATE M23:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=4.54e-06  SB=6.6e-07  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 M24:DRN M24:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=4.28e-06  SB=9.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM25 vdd M25:GATE M25:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=4.04e-06  SB=1.16e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM26 M26:DRN M26:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=3.78e-06  SB=1.42e-06  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM27 vdd M27:GATE M27:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=3.54e-06  SB=1.66e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM28 M28:DRN M28:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.25e-06  SB=1.91e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM29 vdd M29:GATE M29:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.99e-06  SB=2.17e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM40 M40:DRN M40:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=5.04e-06  NRD=2.099  NRS=0.532  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.76e-06  SB=2.44e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.5e-06  SB=2.7e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=5.04e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.24e-06  SB=2.96e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=4.78e-06  SB=4.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.98e-06  SB=3.22e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=4.54e-06  SB=6.6e-07  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.72e-06  SB=3.48e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=4.28e-06  SB=9.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vss M15:GATE M15:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.46e-06  SB=3.74e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=4.04e-06  SB=1.16e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.2e-06  SB=4e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=3.78e-06  SB=1.42e-06  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 vss M17:GATE M17:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.4e-07  SB=4.26e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=3.54e-06  SB=1.66e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M18:DRN M18:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=4.52e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.28e-06  SB=1.92e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vss M19:GATE M19:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=4.78e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.02e-06  SB=2.18e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM30 M30:DRN M30:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.76e-06  SB=2.44e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM31 vdd M31:GATE M31:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.5e-06  SB=2.7e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM32 M32:DRN M32:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.24e-06  SB=2.96e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM33 vdd M33:GATE M33:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.98e-06  SB=3.22e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM34 M34:DRN M34:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.72e-06  SB=3.48e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM35 vdd M35:GATE M35:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.46e-06  SB=3.74e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM36 M36:DRN M36:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.2e-06  SB=4e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM37 vdd M37:GATE M37:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.4e-07  SB=4.26e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM38 M38:DRN M38:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=4.52e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM39 vdd M39:GATE M39:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=4.78e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 ZN ZN:6 0.10123 
R1 ZN:1 ZN:6 0.60627 
R2 M10:DRN ZN:6 15.0394 
R3 ZN:2 ZN:6 0.14337 
R4 M8:DRN ZN:6 25.0255 
R5 M6:DRN ZN:6 50.7459 
R6 ZN:6 M12:DRN 14.9999 
CC13510 ZN:6 I:2 2.21e-18
CC13530 ZN:6 I:6 1.26e-18
CC13776 ZN:6 I 4.44e-18
CC13547 ZN:6 I:9 1.7065e-16
CC13514 ZN:6 I:3 2.26e-18
CC13783 ZN:6 M11:GATE 2.1e-18
CC13526 ZN:6 I:5 1.9005e-16
CC13780 ZN:6 M12:GATE 1.221e-17
CC13721 ZN:6 M18:GATE 1.563e-17
CC13718 ZN:6 M17:GATE 1.406e-17
CC13647 ZN:6 I:18 1.1796e-16
CC13713 ZN:6 M16:GATE 1.566e-17
CC13652 ZN:6 I:19 2.72e-18
CC13712 ZN:6 M15:GATE 1.406e-17
CC13620 ZN:6 I:16 2.51e-18
CC13624 ZN:6 I:17 2.35e-18
CC13724 ZN:6 M19:GATE 1.376e-17
CC13675 ZN:6 M9:GATE 1.307e-17
CC13701 ZN:6 M1:GATE 3.13e-18
CC13677 ZN:6 M8:GATE 1.215e-17
CC13698 ZN:6 M2:GATE 1.21e-17
CC13682 ZN:6 M7:GATE 1.284e-17
CC13695 ZN:6 M3:GATE 1.281e-17
CC13685 ZN:6 M6:GATE 1.29e-17
CC13692 ZN:6 M4:GATE 1.26e-17
CC13687 ZN:6 M5:GATE 1.238e-17
CC13657 ZN:6 I:20 4.89e-18
CC13661 ZN:6 I:21 1.32e-18
CC13667 ZN:6 M20:GATE 4.07e-18
CC13706 ZN:6 M14:GATE 1.566e-17
CC13672 ZN:6 M10:GATE 1.316e-17
CC13703 ZN:6 M13:GATE 1.311e-17
CC13758 ZN:6 M33:GATE 1.32e-18
CC13551 ZN:6 M30:GATE 2.31e-18
CC13768 ZN:6 M31:GATE 6.12e-18
CC13764 ZN:6 M32:GATE 2.11e-18
CC13602 ZN:6 I:12 2.7e-18
CC13606 ZN:6 I:13 6.5e-18
CC13615 ZN:6 I:15 3.34e-18
CC13597 ZN:6 I:11 2.72e-18
R7 M12:DRN M11:SRC 0.001 
CC13778 M12:DRN M12:GATE 1.269e-17
CC13781 M12:DRN M11:GATE 1.975e-17
CC13639 M12:DRN I:18 4.784e-17
CC13761 M12:DRN M32:GATE 3.79e-18
CC13604 M12:DRN I:13 2.362e-17
R8 ZN:1 M6:DRN 21.6929 
R9 M6:DRN M5:SRC 0.001 
CC13522 M6:DRN I:5 1.09e-18
CC13508 M6:DRN I:2 3.761e-17
CC13642 M6:DRN I:18 1.643e-17
CC13684 M6:DRN M6:GATE 8.12e-18
CC13688 M6:DRN M5:GATE 4.57e-18
CC13594 M6:DRN I:11 4.046e-17
R10 ZN:3 ZN:5 0.49643 
R11 ZN ZN:5 0.104 
R12 M28:DRN ZN:5 42.894 
R13 M30:DRN ZN:5 20.8115 
R14 M32:DRN ZN:5 14.9999 
R15 ZN:5 ZN:4 0.22568 
CC13546 ZN:5 I:9 1.2521e-16
CC13775 ZN:5 I 8.14e-18
CC13525 ZN:5 I:5 1.354e-16
CC13646 ZN:5 I:18 5.054e-17
CC13730 ZN:5 M39:GATE 1.65e-17
CC13726 ZN:5 M40:GATE 5.01e-18
CC13762 ZN:5 M32:GATE 1.448e-17
CC13565 ZN:5 M27:GATE 1.799e-17
CC13569 ZN:5 M26:GATE 1.695e-17
CC13757 ZN:5 M33:GATE 1.507e-17
CC13574 ZN:5 M25:GATE 1.799e-17
CC13578 ZN:5 M24:GATE 1.695e-17
CC13753 ZN:5 M34:GATE 1.853e-17
CC13550 ZN:5 M30:GATE 1.649e-17
CC13555 ZN:5 M29:GATE 1.716e-17
CC13767 ZN:5 M31:GATE 1.504e-17
CC13560 ZN:5 M28:GATE 1.724e-17
CC13739 ZN:5 M37:GATE 1.67e-17
CC13735 ZN:5 M38:GATE 1.855e-17
CC13583 ZN:5 M23:GATE 1.792e-17
CC13588 ZN:5 M22:GATE 1.676e-17
CC13748 ZN:5 M35:GATE 1.67e-17
CC13592 ZN:5 M21:GATE 4.38e-18
CC13744 ZN:5 M36:GATE 1.853e-17
R16 M38:DRN ZN:4 15.7136 
R17 M40:DRN ZN:4 15.9027 
R18 M36:DRN ZN:4 15.5311 
R19 ZN:4 M34:DRN 14.9999 
R20 M34:DRN M33:SRC 0.001 
CC13541 M34:DRN I:9 1.59e-18
CC13628 M34:DRN I:18 1.114e-17
CC13755 M34:DRN M33:GATE 4.553e-17
CC13752 M34:DRN M34:GATE 4.557e-17
R21 M36:DRN M35:SRC 0.001 
CC13540 M36:DRN I:9 1.59e-18
CC13627 M36:DRN I:18 1.114e-17
CC13746 M36:DRN M35:GATE 4.495e-17
CC13743 M36:DRN M36:GATE 4.557e-17
R22 M32:DRN M31:SRC 0.001 
CC13629 M32:DRN I:18 1.097e-17
CC13760 M32:DRN M32:GATE 4.497e-17
CC13765 M32:DRN M31:GATE 4.489e-17
R23 ZN:1 M8:DRN 38.3426 
R24 M8:DRN M7:SRC 0.001 
CC13521 M8:DRN I:5 1.09e-18
CC13511 M8:DRN I:3 3.7e-17
CC13641 M8:DRN I:18 1.643e-17
CC13679 M8:DRN M8:GATE 4.57e-18
CC13680 M8:DRN M7:GATE 8.03e-18
CC13613 M8:DRN I:15 4.121e-17
R25 ZN:1 M2:DRN 15.1792 
R26 M2:DRN M1:SRC 0.001 
CC13524 M2:DRN I:5 1.09e-18
CC13504 M2:DRN I:1 4.119e-17
CC13644 M2:DRN I:18 1.614e-17
CC13650 M2:DRN I:19 4.03e-17
CC13700 M2:DRN M2:GATE 4.59e-18
CC13702 M2:DRN M1:GATE 4.8e-18
R27 ZN:3 M30:DRN 54.9921 
R28 M30:DRN M29:SRC 0.001 
CC13515 M30:DRN I:5 1.27e-18
CC13630 M30:DRN I:18 1.111e-17
CC13549 M30:DRN M30:GATE 4.473e-17
CC13553 M30:DRN M29:GATE 4.485e-17
R29 M38:DRN M40:DRN 664.568 
R30 M40:DRN M39:SRC 0.001 
CC13538 M40:DRN I:9 1.56e-18
CC13728 M40:DRN M39:GATE 4.484e-17
CC13625 M40:DRN I:18 1.105e-17
CC13725 M40:DRN M40:GATE 4.595e-17
R31 M38:DRN M37:SRC 0.001 
CC13539 M38:DRN I:9 1.59e-18
CC13626 M38:DRN I:18 1.114e-17
CC13737 M38:DRN M37:GATE 4.495e-17
CC13734 M38:DRN M38:GATE 4.557e-17
R32 M16:DRN ZN:2 15.5479 
R33 M18:DRN ZN:2 15.9319 
R34 M14:DRN ZN:2 14.9999 
R35 ZN:2 M20:SRC 16.1299 
R36 M16:DRN M20:SRC 1298.17 
R37 M18:DRN M20:SRC 645.076 
R38 M20:SRC M19:SRC 0.001 
CC13542 M20:SRC I:9 1.14e-18
CC13535 M20:SRC I:8 2.723e-17
CC13722 M20:SRC M19:GATE 4.59e-18
CC13635 M20:SRC I:18 1.614e-17
CC13662 M20:SRC I:22 4.082e-17
CC13669 M20:SRC M20:GATE 1.913e-17
R39 ZN:1 M4:DRN 14.9999 
R40 M4:DRN M3:SRC 0.001 
CC13523 M4:DRN I:5 1.09e-18
CC13643 M4:DRN I:18 1.643e-17
CC13621 M4:DRN I:17 4.046e-17
CC13696 M4:DRN M3:GATE 4.57e-18
CC13691 M4:DRN M4:GATE 4.57e-18
CC13618 M4:DRN I:16 4.117e-17
R41 M14:DRN M13:SRC 0.001 
CC13545 M14:DRN I:9 1.38e-18
CC13638 M14:DRN I:18 1.643e-17
CC13655 M14:DRN I:20 4.077e-17
CC13708 M14:DRN M14:GATE 4.57e-18
CC13705 M14:DRN M13:GATE 5.3e-18
CC13603 M14:DRN I:13 4.096e-17
R42 ZN:3 M28:DRN 23.447 
R43 M28:DRN M27:SRC 0.001 
CC13516 M28:DRN I:5 1.59e-18
CC13631 M28:DRN I:18 1.114e-17
CC13559 M28:DRN M28:GATE 4.474e-17
CC13563 M28:DRN M27:GATE 4.48e-17
R44 ZN:3 M24:DRN 15.3453 
R45 M22:DRN M24:DRN 1341.25 
R46 M24:DRN M23:SRC 0.001 
CC13518 M24:DRN I:5 1.59e-18
CC13633 M24:DRN I:18 1.114e-17
CC13577 M24:DRN M24:GATE 4.47e-17
CC13581 M24:DRN M23:GATE 4.48e-17
R47 ZN:3 M26:DRN 14.9999 
R48 M26:DRN M25:SRC 0.001 
CC13517 M26:DRN I:5 1.59e-18
CC13632 M26:DRN I:18 1.114e-17
CC13568 M26:DRN M26:GATE 4.47e-17
CC13572 M26:DRN M25:GATE 4.48e-17
R49 ZN:3 M22:DRN 15.5227 
R50 M22:DRN M21:SRC 0.001 
CC13519 M22:DRN I:5 1.53e-18
CC13634 M22:DRN I:18 1.097e-17
CC13587 M22:DRN M22:GATE 4.458e-17
CC13591 M22:DRN M21:GATE 4.593e-17
R51 M10:DRN M9:SRC 0.001 
CC13640 M10:DRN I:18 2.648e-17
CC13671 M10:DRN M10:GATE 8.21e-18
CC13673 M10:DRN M9:GATE 4.93e-18
CC13599 M10:DRN I:12 6.756e-17
R52 M16:DRN M18:DRN 1282.24 
R53 M18:DRN M17:SRC 0.001 
CC13543 M18:DRN I:9 1.38e-18
CC13720 M18:DRN M18:GATE 4.57e-18
CC13716 M18:DRN M17:GATE 4.57e-18
CC13636 M18:DRN I:18 1.643e-17
CC13659 M18:DRN I:21 4.077e-17
CC13607 M18:DRN I:14 4.067e-17
R54 M16:DRN M15:SRC 0.001 
CC13544 M16:DRN I:9 1.38e-18
CC13531 M16:DRN I:7 3.789e-17
CC13528 M16:DRN I:6 3.838e-17
CC13715 M16:DRN M16:GATE 6.96e-18
CC13637 M16:DRN I:18 1.643e-17
CC13709 M16:DRN M15:GATE 7.34e-18
CC13645 ZN I:18 1.86e-18
C55 ZN:6 0 4.8515e-16
C56 M12:DRN 0 4.5e-18
C57 M6:DRN 0 4.5e-18
C58 ZN:5 0 4.8785e-16
C59 M34:DRN 0 7.83e-18
C60 M36:DRN 0 6.46e-18
C61 M32:DRN 0 8.09e-18
C62 M8:DRN 0 4.5e-18
C63 M2:DRN 0 7.52e-18
C64 M30:DRN 0 8.02e-18
C65 M40:DRN 0 9.94e-18
C66 M38:DRN 0 6.66e-18
C67 ZN:2 0 3.6e-19
C68 M20:SRC 0 7.29e-18
C69 M4:DRN 0 4.5e-18
C70 M14:DRN 0 4.85e-18
C71 M28:DRN 0 6.34e-18
C72 M24:DRN 0 6.61e-18
C73 M26:DRN 0 6.43e-18
C74 M22:DRN 0 1.074e-17
C75 M10:DRN 0 5.2e-18
C76 ZN:1 0 3.4e-19
C77 M18:DRN 0 4.5e-18
C78 M16:DRN 0 4.5e-18
C79 ZN 0 5.7e-19
R80 M3:GATE I:17 86.5669 
R81 M23:GATE I:17 111.3 
R82 I:1 I:17 2249.74 
R83 I:4 I:17 22.6743 
R84 I:16 I:17 21.5119 
R85 I:17 I:19 20.8471 
R86 I:1 I:19 22.0055 
R87 I:4 I:19 23.1435 
R88 M2:GATE I:19 85.0652 
R89 I:19 M22:GATE 111.3 
R90 M19:GATE I:22 83.8364 
R91 M39:GATE I:22 101.061 
R92 I:8 I:22 22.3658 
R93 I:21 I:22 21.5119 
R94 I:10 I:22 32.926 
R95 I:22 I 68.4613 
R96 I:8 I 34.0542 
R97 I I:10 0.70947 
R98 I:9 I:10 0.69247 
R99 I:8 I:10 64.0913 
R100 I:21 I:10 22 
R101 I:14 I:10 29.8079 
R102 I:10 I:6 118.673 
R103 I:9 I:6 29.3535 
R104 I:7 I:6 31.0275 
R105 M16:GATE I:6 94.0755 
R106 M36:GATE I:6 111.3 
R107 I:6 I:14 33.904 
R108 M17:GATE I:14 82.8124 
R109 I:9 I:14 45.4767 
R110 M37:GATE I:14 100.037 
R111 I:14 I:21 21.9794 
R112 M38:GATE I:21 103.792 
R113 I:21 M18:GATE 86.5669 
R114 M40:GATE I:8 97.7846 
R115 I:8 M20:GATE 80.5597 
R116 M29:GATE I:12 111.3 
R117 M9:GATE I:12 85.0652 
R118 M10:GATE I:12 222.334 
R119 M30:GATE I:12 263.044 
R120 I:5 I:12 23.3308 
R121 I:18 I:12 57.4715 
R122 I:12 I:15 21.9469 
R123 M28:GATE I:15 111.3 
R124 I:5 I:15 18.0836 
R125 I:3 I:15 35.539 
R126 I:15 M8:GATE 81.2035 
R127 M12:GATE M32:GATE 1092.88 
R128 I:13 M32:GATE 266.204 
R129 M32:GATE I:18 282.501 
R130 M12:GATE I:18 238.78 
R131 M31:GATE I:18 88.7752 
R132 M10:GATE I:18 240.862 
R133 M30:GATE I:18 284.964 
R134 I:13 I:18 58.1624 
R135 I:18 M11:GATE 94.0755 
R136 M13:GATE I:13 86.5669 
R137 I:9 I:13 23.3292 
R138 I:7 I:13 4229.71 
R139 M33:GATE I:13 103.792 
R140 M12:GATE I:13 225.005 
R141 I:13 I:20 21.9521 
R142 M34:GATE I:20 99.1711 
R143 I:9 I:20 18.3541 
R144 I:7 I:20 34.7786 
R145 I:20 M14:GATE 81.9458 
R146 M7:GATE I:3 94.0755 
R147 M27:GATE I:3 111.3 
R148 I:2 I:3 28.1628 
R149 I:3 I:5 24.3077 
R150 I:4 I:5 0.69451 
R151 I:2 I:5 29.9639 
R152 I:5 I:11 44.302 
R153 M25:GATE I:11 111.3 
R154 M5:GATE I:11 81.9458 
R155 I:4 I:11 29.5529 
R156 I:2 I:11 34.9924 
R157 I:11 I:16 21.5119 
R158 M24:GATE I:16 111.3 
R159 I:4 I:16 22 
R160 I:16 M4:GATE 83.8364 
R161 M6:GATE I:2 94.0755 
R162 M26:GATE I:2 111.3 
R163 I:2 I:4 125.543 
R164 I:4 I:1 23.3838 
R165 M21:GATE I:1 111.3 
R166 I:1 M1:GATE 81.2035 
R167 M30:GATE M10:GATE 1102.4 
R168 M15:GATE I:7 94.0755 
R169 M35:GATE I:7 111.3 
R170 I:7 I:9 23.7964 
C171 M3:GATE 0 2.388e-17
C172 I:17 0 2.47e-18
C173 I:19 0 2.8e-18
C174 M22:GATE 0 3.824e-17
C175 M19:GATE 0 3.121e-17
C176 I:22 0 4.14e-18
C177 I 0 6.732e-17
C178 I:10 0 1.27e-17
C179 I:6 0 2.92e-18
C180 I:14 0 4.57e-18
C181 I:21 0 4.46e-18
C182 M18:GATE 0 2.854e-17
C183 M40:GATE 0 6.44e-17
C184 I:8 0 3.337e-17
C185 M20:GATE 0 2.789e-17
C186 M29:GATE 0 1.486e-17
C187 I:12 0 5.08e-18
C188 I:15 0 1.161e-17
C189 M8:GATE 0 2.869e-17
C190 M37:GATE 0 3.47e-17
C191 M32:GATE 0 3.365e-17
C192 I:18 0 1.715e-16
C193 M11:GATE 0 2.716e-17
C194 M36:GATE 0 3.237e-17
C195 M39:GATE 0 3.91e-17
C196 M2:GATE 0 3.319e-17
C197 M16:GATE 0 1.978e-17
C198 M13:GATE 0 2.222e-17
C199 I:13 0 4.58e-18
C200 I:20 0 9.18e-18
C201 M14:GATE 0 2.583e-17
C202 M7:GATE 0 2.318e-17
C203 I:3 0 4.26e-18
C204 I:5 0 3.526e-17
C205 I:11 0 2.83e-18
C206 I:16 0 2.73e-18
C207 M4:GATE 0 2.886e-17
C208 M6:GATE 0 2.261e-17
C209 I:2 0 2.19e-18
C210 I:4 0 2.052e-17
C211 I:1 0 2.661e-17
C212 M1:GATE 0 5.066e-17
C213 M30:GATE 0 1.664e-17
C214 M10:GATE 0 2.655e-17
C215 M31:GATE 0 3.67e-17
C216 M38:GATE 0 4.118e-17
C217 M28:GATE 0 1.484e-17
C218 M5:GATE 0 2.262e-17
C219 M12:GATE 0 2.313e-17
C220 M33:GATE 0 3.139e-17
C221 M15:GATE 0 2.343e-17
C222 I:7 0 4.33e-18
C223 I:9 0 1.243e-17
C224 M9:GATE 0 2.207e-17
C225 M35:GATE 0 3.513e-17
C226 M34:GATE 0 3.927e-17
C227 M24:GATE 0 3.54e-17
C228 M25:GATE 0 2.887e-17
C229 M21:GATE 0 7.888e-17
C230 M23:GATE 0 3.081e-17
C231 M27:GATE 0 2.919e-17
C232 M17:GATE 0 2.296e-17
C233 M26:GATE 0 2.945e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
