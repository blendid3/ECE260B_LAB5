.SUBCKT NR2D2 A1 A2 ZN
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.93e-07  AD=7.4e-14  AS=3.9e-14  PD=1.16e-06  PS=5.9e-07  SA=9.7e-07  SB=1.9e-07  NRD=0.619  NRS=4.183  SCA=11.516  SCB=0.012  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.1e-07  SB=4.5e-07  NRD=4.183  NRS=4.183  SCA=11.516  SCB=0.012  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.5e-07  SB=7.1e-07  NRD=4.183  NRS=4.183  SCA=11.516  SCB=0.012  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.93e-07  AD=3.9e-14  AS=7.4e-14  PD=5.9e-07  PS=1.16e-06  SA=1.9e-07  SB=9.7e-07  NRD=4.183  NRS=0.619  SCA=11.516  SCB=0.012  SCC=0.001 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=5.3e-07  AD=1.11e-13  AS=5.3e-14  PD=1.48e-06  PS=7.3e-07  SA=9.9e-07  SB=2.1e-07  NRD=0.571  NRS=1.971  SCA=9.514  SCB=0.01  SCC=0.0008075 
MMM6 M5:SRC M6:GATE M6:SRC vdd pch L=6e-08 W=5.3e-07  AD=5.3e-14  AS=5.3e-14  PD=7.3e-07  PS=7.3e-07  SA=7.3e-07  SB=4.7e-07  NRD=1.971  NRS=2.063  SCA=9.514  SCB=0.01  SCC=0.0008075 
MMM7 M7:DRN M7:GATE M7:SRC vdd pch L=6e-08 W=5.3e-07  AD=5.3e-14  AS=5.3e-14  PD=7.3e-07  PS=7.3e-07  SA=4.7e-07  SB=7.3e-07  NRD=2.063  NRS=1.971  SCA=9.514  SCB=0.01  SCC=0.0008075 
MMM8 M7:SRC M8:GATE vdd vdd pch L=6e-08 W=5.3e-07  AD=5.3e-14  AS=1.11e-13  PD=7.3e-07  PS=1.48e-06  SA=2.1e-07  SB=9.9e-07  NRD=1.971  NRS=0.571  SCA=9.514  SCB=0.01  SCC=0.0008075 
R0 M2:DRN M1:SRC 0.001 
R1 M3:SRC M1:SRC 2653.91 
R2 M1:SRC ZN 31.5288 
CC47660 M1:SRC M2:GATE 2.824e-17
CC47630 M1:SRC M1:GATE 1.03e-18
CC47631 M1:SRC A2 3.052e-17
R3 M6:SRC ZN 30.8733 
R4 ZN M3:SRC 30.959 
CC47657 ZN A1 7.755e-17
CC47639 ZN A1:1 9.64e-18
CC47662 ZN M2:GATE 6.61e-18
CC47650 ZN M6:GATE 3.66e-18
CC47644 ZN M7:GATE 8e-18
CC47667 ZN M3:GATE 5.32e-18
CC47624 ZN M8:GATE 4.68e-18
CC47625 ZN M4:GATE 7.39e-18
CC47626 ZN M1:GATE 2.83e-18
CC47627 ZN A2 1.5663e-16
R5 M3:SRC M4:DRN 0.001 
CC47636 M3:SRC A1:1 2.731e-17
CC47665 M3:SRC M3:GATE 1.07e-18
CC47628 M3:SRC M4:GATE 1.024e-17
CC47629 M3:SRC A2 2.032e-17
R6 M6:SRC M7:DRN 0.001 
CC47634 M6:SRC A1:1 8.52e-18
CC47642 M6:SRC M7:GATE 2.769e-17
CC47652 M6:SRC A1 3.03e-18
CC47647 M6:SRC M6:GATE 2.806e-17
CC47622 M6:SRC M5:GATE 1.04e-18
CC47623 M6:SRC A2 5.02e-18
C7 M1:SRC 0 8.27e-18
C8 ZN 0 1.1149e-16
C9 M3:SRC 0 7.54e-18
C10 M6:SRC 0 6.52e-18
R11 A2 M8:GATE 147.192 
R12 M8:GATE M4:GATE 535.777 
CC47641 M8:GATE M7:GATE 1.317e-17
CC47633 M8:GATE A1:1 9.07e-18
R13 M4:GATE A2 121.333 
CC47635 M4:GATE A1:1 2.2e-18
CC47664 M4:GATE M3:GATE 4.58e-18
R14 M1:GATE A2 125.984 
R15 A2 M5:GATE 152.833 
CC47645 A2 M7:GATE 9.67e-18
CC47640 A2 A1:1 3.69e-18
CC47663 A2 M2:GATE 2.54e-18
CC47651 A2 M6:GATE 9.71e-18
CC47658 A2 A1 2.258e-17
R16 M5:GATE M1:GATE 499.026 
CC47648 M5:GATE M6:GATE 1.33e-17
CC47649 M1:GATE M6:GATE 5.17e-18
CC47638 M1:GATE A1:1 8.67e-18
CC47661 M1:GATE M2:GATE 3.11e-18
C17 M8:GATE 0 7.313e-17
C18 M4:GATE 0 4.352e-17
C19 A2 0 2.6477e-16
C20 M5:GATE 0 8.65e-17
C21 M1:GATE 0 5.106e-17
R22 M3:GATE A1:1 95.3999 
R23 M7:GATE A1:1 112.625 
R24 M6:GATE A1:1 242.549 
R25 M2:GATE A1:1 205.452 
R26 A1:1 A1 38.351 
R27 M6:GATE A1 438.864 
R28 A1 M2:GATE 371.746 
R29 M2:GATE M6:GATE 745.524 
C30 A1:1 0 4.721e-17
C31 A1 0 1.615e-17
C32 M2:GATE 0 3.262e-17
C33 M6:GATE 0 3.976e-17
C34 M7:GATE 0 4.039e-17
C35 M3:GATE 0 5.423e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
