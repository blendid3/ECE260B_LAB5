.SUBCKT OR2D4 A1 A2 Z
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.3e-14  PD=7.2e-07  PS=7.25e-07  SA=1.75e-06  SB=4.2e-07  NRD=2.057  NRS=1.092  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.3e-14  AS=5.2e-14  PD=7.25e-07  PS=7.2e-07  SA=1.485e-06  SB=6.85e-07  NRD=1.092  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.266e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.5e-14  PD=7.2e-07  PS=7.3e-07  SA=1.225e-06  SB=9.45e-07  NRD=2.057  NRS=0.702  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4e-14  PD=5.9e-07  PS=5.95e-07  SA=9.62e-07  SB=4.2e-07  NRD=4.141  NRS=3.415  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.5e-14  AS=5.1e-14  PD=7.3e-07  PS=7.15e-07  SA=9.55e-07  SB=1.215e-06  NRD=0.702  NRS=3.014  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=4e-14  AS=3.9e-14  PD=5.95e-07  PS=5.9e-07  SA=6.3e-07  SB=6.85e-07  NRD=3.415  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M13:SRC M14:GATE M14:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.1e-14  AS=5.3e-14  PD=7.15e-07  PS=7.25e-07  SA=7e-07  SB=1.47e-06  NRD=3.014  NRS=1.092  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=4e-14  PD=5.9e-07  PS=7.6e-07  SA=2.54e-07  SB=9.45e-07  NRD=4.141  NRS=11.621  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 M14:SRC M15:GATE M15:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.3e-14  AS=5.2e-14  PD=7.25e-07  PS=7.2e-07  SA=4.35e-07  SB=1.735e-06  NRD=1.092  NRS=2.009  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=2.09e-07  AD=2e-14  AS=2e-14  PD=3.8e-07  PS=4.05e-07  SA=1.005e-06  SB=1.185e-06  NRD=0.694  NRS=5.196  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM16 M15:SRC M16:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=9.1e-14  PD=7.2e-07  PS=1.39e-06  SA=1.75e-07  SB=1.995e-06  NRD=2.099  NRS=0.541  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M5:SRC M6:GATE vss vss nch L=6e-08 W=1.95e-07  AD=2e-14  AS=2.3e-14  PD=4.05e-07  PS=4.35e-07  SA=7.35e-07  SB=1.455e-06  NRD=5.196  NRS=0.634  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=1.95e-07  AD=2.3e-14  AS=2e-14  PD=4.35e-07  PS=3.95e-07  SA=4.35e-07  SB=1.755e-06  NRD=0.634  NRS=8.262  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM8 M7:SRC M8:GATE vss vss nch L=6e-08 W=1.95e-07  AD=2e-14  AS=3.4e-14  PD=3.95e-07  PS=7.4e-07  SA=1.75e-07  SB=2.015e-06  NRD=8.262  NRS=0.947  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=2.01e-06  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M11:SRC M12:DRN 0.001 
R1 M10:DRN M12:DRN 1622.9 
R2 M12:DRN Z 15.7158 
CC11745 M12:DRN A2 1.32e-18
CC11754 M12:DRN N_13:1 1.581e-17
CC11775 M12:DRN M11:GATE 4.786e-17
CC11771 M12:DRN M12:GATE 4.642e-17
R3 M4:DRN Z 15.6351 
R4 M10:DRN Z 15.362 
R5 Z M2:DRN 15.2927 
CC11744 Z M13:GATE 1.32e-18
CC11747 Z A2 2.508e-17
CC11798 Z M7:SRC 2.729e-17
CC11794 Z M4:GATE 1.62e-18
CC11791 Z M3:GATE 4.23e-18
CC11787 Z M1:GATE 3.46e-18
CC11785 Z M2:GATE 2.17e-18
CC11784 Z M9:GATE 6.01e-18
CC11766 Z N_13:2 8.78e-18
CC11760 Z N_13:1 8.806e-17
CC11749 Z M5:GATE 1.29e-18
CC11780 Z M10:GATE 8.16e-18
CC11778 Z M11:GATE 1.014e-17
CC11772 Z M12:GATE 5.29e-18
R6 M2:DRN M1:SRC 0.001 
CC11788 M2:DRN M1:GATE 1.834e-17
CC11786 M2:DRN M2:GATE 4.182e-17
CC11765 M2:DRN N_13:2 3.993e-17
CC11759 M2:DRN N_13:1 1.495e-17
R7 M10:DRN M9:SRC 0.001 
CC11783 M10:DRN M9:GATE 4.599e-17
CC11782 M10:DRN M10:GATE 4.742e-17
CC11763 M10:DRN N_13:2 1.66e-18
CC11755 M10:DRN N_13:1 1.302e-17
R8 M4:DRN M3:SRC 0.001 
CC11793 M4:DRN M4:GATE 8.27e-18
CC11790 M4:DRN M3:GATE 8.56e-18
CC11764 M4:DRN N_13:2 1.633e-17
CC11758 M4:DRN N_13:1 8.494e-17
C9 M12:DRN 0 1.122e-17
C10 Z 0 2.9243e-16
C11 M2:DRN 0 1.008e-17
C12 M10:DRN 0 9.22e-18
C13 M4:DRN 0 1.005e-17
CC11751 M13:SRC A2 1.08e-18
R14 A2 M16:GATE 141.439 
R15 M16:GATE M8:GATE 692.091 
CC11812 M16:GATE M15:GATE 1.352e-17
CC11802 M16:GATE A1:1 9.13e-18
CC11752 M16:GATE N_13:1 5.38e-18
R16 M8:GATE A2 153.531 
CC11835 M8:GATE M7:GATE 1.36e-18
CC11808 M8:GATE A1:1 8.54e-18
CC11797 M8:GATE M7:SRC 2.43e-17
R17 M5:GATE A2 157.725 
R18 A2 M13:GATE 145.139 
CC11833 A2 M6:GATE 7.88e-18
CC11827 A2 A1 3.02e-17
CC11820 A2 M14:GATE 1.15e-18
CC11815 A2 M15:GATE 1.074e-17
CC11810 A2 A1:1 1.685e-17
CC11801 A2 M5:SRC 1.3362e-16
CC11799 A2 M7:SRC 6.751e-17
CC11795 A2 M4:GATE 4.21e-18
CC11773 A2 M12:GATE 7.67e-18
CC11769 A2 M14:SRC 5.43e-18
CC11761 A2 N_13:1 1.339e-17
R19 M13:GATE M5:GATE 625.41 
CC11818 M13:GATE M14:GATE 3.28e-18
CC11806 M13:GATE A1:1 1.859e-17
CC11753 M13:GATE N_13:1 7.97e-18
CC11770 M13:GATE M12:GATE 1.1e-17
CC11768 M13:GATE M14:SRC 3.76e-18
CC11831 M5:GATE M6:GATE 1.12e-18
CC11757 M5:GATE N_13:1 1.035e-17
CC11800 M5:GATE M5:SRC 2.445e-17
CC11792 M5:GATE M4:GATE 2.87e-18
C20 M16:GATE 0 7.913e-17
C21 M8:GATE 0 4.429e-17
C22 A2 0 2.059e-16
C23 M13:GATE 0 5.768e-17
C24 M5:GATE 0 3.458e-17
R25 M4:GATE N_13:1 80.5597 
R26 M14:SRC N_13:1 102.139 
R27 M5:SRC N_13:1 98.3435 
R28 M7:SRC N_13:1 100.431 
R29 M3:GATE N_13:1 207.507 
R30 M11:GATE N_13:1 245.499 
R31 M12:GATE N_13:1 111.3 
R32 N_13:1 N_13:2 54.6703 
CC11821 N_13:1 M14:GATE 6.94e-18
CC11816 N_13:1 M15:GATE 2.35e-18
CC11839 N_13:1 M7:GATE 2.44e-18
R33 M2:GATE N_13:2 94.0755 
R34 M10:GATE N_13:2 111.3 
R35 M3:GATE N_13:2 255.763 
R36 M11:GATE N_13:2 302.591 
R37 M9:GATE N_13:2 164.389 
R38 N_13:2 M1:GATE 138.947 
R39 M1:GATE M9:GATE 635.948 
R40 M11:GATE M3:GATE 1148.51 
R41 M14:SRC M7:SRC 136.128 
R42 M7:SRC M5:SRC 131.069 
CC11836 M7:SRC M7:GATE 2.623e-17
CC11809 M7:SRC A1:1 1.738e-17
CC11825 M7:SRC A1 1.085e-17
R43 M5:SRC M14:SRC 133.299 
CC11830 M5:SRC M6:GATE 2.443e-17
CC11826 M5:SRC A1 4.46e-18
CC11804 M14:SRC A1:1 3.994e-17
CC11823 M14:SRC A1 8.085e-17
CC11813 M14:SRC M15:GATE 2.586e-17
C44 N_13:1 0 9.994e-17
C45 N_13:2 0 6.184e-17
C46 M1:GATE 0 6.417e-17
C47 M9:GATE 0 1.0192e-16
C48 M12:GATE 0 4.67e-17
C49 M11:GATE 0 7.971e-17
C50 M3:GATE 0 6.471e-17
C51 M10:GATE 0 7.134e-17
C52 M7:SRC 0 2.273e-17
C53 M5:SRC 0 5.22e-18
C54 M14:SRC 0 3.786e-17
C55 M4:GATE 0 3.683e-17
C56 M2:GATE 0 2.364e-17
R57 M7:GATE A1:1 119.78 
R58 M15:GATE A1:1 111.3 
R59 M14:GATE A1:1 210.63 
R60 M6:GATE A1:1 226.678 
R61 A1:1 A1 33.6214 
R62 M14:GATE A1 521.52 
R63 A1 M6:GATE 561.257 
R64 M6:GATE M14:GATE 895.065 
C65 A1:1 0 3.053e-17
C66 A1 0 7.52e-18
C67 M6:GATE 0 4.083e-17
C68 M14:GATE 0 5.229e-17
C69 M15:GATE 0 4.117e-17
C70 M7:GATE 0 3.415e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
