.SUBCKT BUFFD8 I Z
MMM20 vdd M20:GATE M20:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.95e-07  SB=2.255e-06  NRD=2.099  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 M20:SRC M21:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.35e-07  SB=2.515e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=9.1e-14  AS=5.2e-14  PD=1.39e-06  PS=7.2e-07  SA=1.75e-07  SB=2.775e-06  NRD=0.541  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M9:SRC M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.35e-07  SB=2.515e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 M11:DRN M11:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.8e-14  AS=3.9e-14  PD=1.13e-06  PS=5.9e-07  SA=1.75e-07  SB=2.775e-06  NRD=0.592  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.97e-07  AD=6.8e-14  AS=3.9e-14  PD=1.13e-06  PS=5.9e-07  SA=2.775e-06  SB=1.75e-07  NRD=0.496  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 vdd M12:GATE M12:SRC vdd pch L=6e-08 W=5.24e-07  AD=9.1e-14  AS=5.2e-14  PD=1.39e-06  PS=7.2e-07  SA=2.775e-06  SB=1.75e-07  NRD=0.446  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.515e-06  SB=4.35e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 M13:DRN M13:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.515e-06  SB=4.35e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.255e-06  SB=6.95e-07  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 vdd M14:GATE M14:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.255e-06  SB=6.95e-07  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.995e-06  SB=9.55e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 M15:DRN M15:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.995e-06  SB=9.55e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.735e-06  SB=1.215e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 vdd M16:GATE M16:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.735e-06  SB=1.215e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.475e-06  SB=1.475e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 M17:DRN M17:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.475e-06  SB=1.475e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.215e-06  SB=1.735e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 vdd M18:GATE M18:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.215e-06  SB=1.735e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.55e-07  SB=1.995e-06  NRD=4.141  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 M19:DRN M19:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.55e-07  SB=1.995e-06  NRD=2.057  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.95e-07  SB=2.255e-06  NRD=4.183  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
R0 M3:SRC Z:2 14.9999 
R1 M6:DRN Z:2 14.9999 
R2 M8:DRN Z:2 15.2796 
R3 Z Z:2 0.03813 
R4 Z:2 M2:DRN 15.2796 
CC78215 Z:2 M9:SRC 2.27e-18
CC78206 Z:2 M2:GATE 9.94e-18
CC78203 Z:2 M3:GATE 1.356e-17
CC78097 Z:2 N_14:2 3.73e-18
CC78162 Z:2 M7:GATE 1.416e-17
CC78157 Z:2 M6:GATE 1.666e-17
CC78152 Z:2 M5:GATE 1.27e-17
CC78138 Z:2 N_14:6 6.075e-17
CC78148 Z:2 M4:GATE 1.489e-17
CC78145 Z:2 M8:GATE 1.9e-18
CC78141 Z:2 M1:GATE 5.92e-18
CC78121 Z:2 N_14:5 5.96e-17
CC78174 Z:2 M18:GATE 1.14e-18
CC78167 Z:2 M19:GATE 1.8e-18
R5 M2:DRN M1:SRC 0.001 
CC78207 M2:DRN M2:GATE 5.07e-18
CC78134 M2:DRN N_14:6 1.0001e-16
CC78140 M2:DRN M1:GATE 5.06e-18
R6 M14:SRC Z:1 14.9999 
R7 M17:DRN Z:1 14.9999 
R8 M19:DRN Z:1 15.2709 
R9 M13:DRN Z:1 15.2709 
R10 Z:1 Z 0.104 
CC78092 Z:1 N_14:1 4.29e-18
CC78098 Z:1 N_14:2 1.9e-18
CC78158 Z:1 M6:GATE 1.43e-18
CC78149 Z:1 M4:GATE 1.03e-18
CC78139 Z:1 N_14:6 9.277e-17
CC78190 Z:1 M13:GATE 1.997e-17
CC78187 Z:1 M14:GATE 1.931e-17
CC78184 Z:1 M15:GATE 2.608e-17
CC78122 Z:1 N_14:5 6.488e-17
CC78181 Z:1 M16:GATE 2.194e-17
CC78178 Z:1 M17:GATE 1.886e-17
CC78124 Z:1 M12:GATE 4.42e-18
CC78175 Z:1 M18:GATE 1.804e-17
CC78168 Z:1 M19:GATE 4.54e-18
R11 M13:DRN M12:SRC 0.001 
CC78189 M13:DRN M13:GATE 4.471e-17
CC78123 M13:DRN M12:GATE 4.583e-17
CC78130 M13:DRN N_14:6 1.38e-17
R12 M8:DRN M7:SRC 0.001 
CC78103 M8:DRN N_14:4 3.491e-17
CC78099 M8:DRN N_14:3 1.785e-17
CC78117 M8:DRN N_14:5 1.63e-18
CC78131 M8:DRN N_14:6 1.387e-17
CC78160 M8:DRN M7:GATE 5.07e-18
CC78144 M8:DRN M8:GATE 3.835e-17
R13 M19:DRN M18:SRC 0.001 
CC78110 M19:DRN N_14:5 1.52e-18
CC78165 M19:DRN M19:GATE 4.577e-17
CC78170 M19:DRN M18:GATE 4.488e-17
CC78127 M19:DRN N_14:6 1.266e-17
R14 M17:DRN M16:SRC 0.001 
CC78179 M17:DRN M16:GATE 4.48e-17
CC78177 M17:DRN M17:GATE 4.531e-17
CC78128 M17:DRN N_14:6 1.265e-17
R15 M14:SRC M15:DRN 0.001 
CC78185 M14:SRC M14:GATE 4.485e-17
CC78183 M14:SRC M15:GATE 4.476e-17
CC78129 M14:SRC N_14:6 1.262e-17
R16 M6:DRN M5:SRC 0.001 
CC78100 M6:DRN N_14:3 2.812e-17
CC78088 M6:DRN N_14:1 5.644e-17
CC78132 M6:DRN N_14:6 1.398e-17
CC78155 M6:DRN M6:GATE 5.69e-18
CC78150 M6:DRN M5:GATE 5.07e-18
R17 M3:SRC M4:DRN 0.001 
CC78205 M3:SRC M3:GATE 5.07e-18
CC78089 M3:SRC N_14:1 2.108e-17
CC78095 M3:SRC N_14:2 6.214e-17
CC78133 M3:SRC N_14:6 1.43e-17
CC78147 M3:SRC M4:GATE 6.92e-18
C18 Z:2 0 1.9451e-16
C19 M2:DRN 0 1.177e-17
C20 Z:1 0 2.1524e-16
C21 Z 0 2.3e-19
C22 M13:DRN 0 1.812e-17
C23 M8:DRN 0 5.28e-18
C24 M19:DRN 0 1.355e-17
C25 M17:DRN 0 4.29e-18
C26 M14:SRC 0 4.29e-18
C27 M6:DRN 0 4.6e-18
C28 M3:SRC 0 4.6e-18
R29 M10:GATE I:1 94.0755 
R30 M9:GATE I:1 193.745 
R31 M20:GATE I:1 229.22 
R32 I I:1 18.0879 
R33 M22:GATE I:1 230.123 
R34 M11:GATE I:1 194.508 
R35 I:1 M21:GATE 111.3 
CC78199 I:1 M20:SRC 1.651e-17
CC78202 I:1 M11:DRN 2.776e-17
CC78214 I:1 M9:SRC 6.896e-17
CC78196 M21:GATE M20:SRC 4.587e-17
CC78108 M21:GATE N_14:5 1.141e-17
R36 I M11:GATE 419.96 
R37 M11:GATE M22:GATE 702.529 
CC78114 M11:GATE N_14:5 7.82e-18
R38 M22:GATE I 496.855 
CC78191 M22:GATE M22:DRN 2.764e-17
CC78107 M22:GATE N_14:5 1.975e-17
CC78125 M22:GATE N_14:6 5.41e-18
R39 M9:GATE I 423.884 
R40 I M20:GATE 501.498 
CC78198 I M20:SRC 1.22e-18
CC78201 I M11:DRN 2.01e-18
CC78213 I M9:SRC 2.998e-17
CC78193 I M22:DRN 1.96e-18
CC78119 I N_14:5 1.199e-16
R41 M20:GATE M9:GATE 702.129 
CC78164 M20:GATE M19:GATE 6.8e-18
CC78197 M20:GATE M20:SRC 4.565e-17
CC78109 M20:GATE N_14:5 7.44e-18
CC78143 M9:GATE M8:GATE 1.1e-18
CC78211 M9:GATE M9:SRC 5.07e-18
CC78116 M9:GATE N_14:5 6.62e-18
CC78102 M9:GATE N_14:4 7.03e-18
CC78210 M10:GATE M9:SRC 5.98e-18
CC78115 M10:GATE N_14:5 7.38e-18
C42 I:1 0 1.507e-17
C43 M21:GATE 0 4.177e-17
C44 M11:GATE 0 5.304e-17
C45 M22:GATE 0 3.39e-17
C46 I 0 2.243e-17
C47 M20:GATE 0 8.373e-17
C48 M9:GATE 0 6.029e-17
C49 M10:GATE 0 3.527e-17
R50 N_14:4 M19:GATE 138.86 
R51 M19:GATE M8:GATE 867.874 
R52 M8:GATE N_14:4 130.181 
R53 N_14:3 N_14:4 22.2465 
R54 M7:GATE N_14:4 184.482 
R55 M18:GATE N_14:4 196.781 
R56 N_14:4 N_14:5 22.6494 
R57 M22:DRN N_14:5 32.9016 
R58 M20:SRC N_14:5 16.0124 
R59 N_14:3 N_14:5 22.8844 
R60 M11:DRN N_14:5 32.3885 
R61 N_14:5 M9:SRC 15.9173 
R62 M9:SRC M11:DRN 907.484 
R63 N_14:3 M18:GATE 284.238 
R64 M18:GATE M7:GATE 2323.11 
R65 M7:GATE N_14:3 266.473 
R66 M6:GATE N_14:3 172.62 
R67 M17:GATE N_14:3 184.128 
R68 N_14:3 N_14:1 42.241 
R69 M5:GATE N_14:1 99.3746 
R70 M16:GATE N_14:1 106 
R71 M6:GATE N_14:1 345.24 
R72 M17:GATE N_14:1 368.257 
R73 N_14:2 N_14:1 60.1649 
R74 M15:GATE N_14:1 262.256 
R75 N_14:1 M4:GATE 245.865 
R76 N_14:2 M4:GATE 245.865 
R77 M4:GATE M15:GATE 1071.73 
R78 M15:GATE N_14:2 262.256 
R79 M3:GATE N_14:2 99.3746 
R80 M14:GATE N_14:2 106 
R81 N_14:2 N_14:6 22.4472 
R82 M2:GATE N_14:6 90.365 
R83 M13:GATE N_14:6 83.475 
R84 M12:GATE N_14:6 139.136 
R85 N_14:6 M1:GATE 113.545 
R86 M1:GATE M12:GATE 808.302 
R87 M17:GATE M6:GATE 1504.89 
R88 M20:SRC M22:DRN 673.372 
C89 M19:GATE 0 4.322e-17
C90 M8:GATE 0 2.69e-17
C91 N_14:4 0 2.671e-17
C92 N_14:5 0 2.0981e-16
C93 M9:SRC 0 9e-18
C94 M11:DRN 0 1.455e-17
C95 M18:GATE 0 4.127e-17
C96 M7:GATE 0 3.285e-17
C97 N_14:3 0 2.2e-19
C98 N_14:1 0 2.33e-18
C99 M4:GATE 0 3.04e-17
C100 M15:GATE 0 3.879e-17
C101 N_14:2 0 1.27e-18
C102 N_14:6 0 1.2213e-16
C103 M1:GATE 0 6.452e-17
C104 M12:GATE 0 8.957e-17
C105 M17:GATE 0 5.039e-17
C106 M6:GATE 0 3.718e-17
C107 M16:GATE 0 4.175e-17
C108 M14:GATE 0 4.17e-17
C109 M13:GATE 0 4.218e-17
C110 M20:SRC 0 1.375e-17
C111 M22:DRN 0 1.897e-17
C112 M3:GATE 0 3.329e-17
C113 M5:GATE 0 3.256e-17
C114 M2:GATE 0 3.463e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
