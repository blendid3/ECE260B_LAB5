.SUBCKT INVD8 I ZN
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.75e-06  SB=4.5e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.49e-06  SB=7.1e-07  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7.4e-14  AS=3.9e-14  PD=1.16e-06  PS=5.9e-07  SA=2.01e-06  SB=1.9e-07  NRD=0.531  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.23e-06  SB=9.7e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.75e-06  SB=4.5e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.7e-07  SB=1.23e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.49e-06  SB=7.1e-07  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7.1e-07  SB=1.49e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.23e-06  SB=9.7e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vdd M15:GATE M15:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.5e-07  SB=1.75e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.7e-07  SB=1.23e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=9.9e-14  PD=7.2e-07  PS=1.42e-06  SA=1.9e-07  SB=2.01e-06  NRD=2.057  NRS=0.554  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7.1e-07  SB=1.49e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.5e-07  SB=1.75e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=7.4e-14  PD=5.9e-07  PS=1.16e-06  SA=1.9e-07  SB=2.01e-06  NRD=4.141  NRS=0.619  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.2e-07  AD=9.9e-14  AS=5.2e-14  PD=1.42e-06  PS=7.2e-07  SA=2.01e-06  SB=1.9e-07  NRD=0.466  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M12:GATE I:1 111.3 
R1 M3:GATE I:1 234.865 
R2 M11:GATE I:1 277.87 
R3 M4:GATE I:1 94.0755 
R4 M13:GATE I:1 273.588 
R5 M5:GATE I:1 231.246 
R6 I:5 I:1 60.9247 
R7 I:1 I:2 59.5436 
CC38383 I:1 M6:DRN 1.552e-17
CC38390 I:1 M4:DRN 6.121e-17
CC38334 I:1 ZN:2 7.36e-18
CC38359 I:1 M12:DRN 1.61e-18
CC38353 I:1 M14:DRN 1.68e-18
R8 M2:GATE I:2 86.5669 
R9 M3:GATE I:2 230.351 
R10 M11:GATE I:2 272.525 
R11 M10:GATE I:2 111.3 
R12 M9:GATE I:2 145.434 
R13 I:2 M1:GATE 107.078 
CC38365 I:2 M10:DRN 4.52e-18
CC38396 I:2 M2:DRN 8.334e-17
CC38391 I:2 M4:DRN 1.678e-17
CC38335 I:2 ZN:2 5.013e-17
CC38360 I:2 M12:DRN 1.63e-18
R14 M1:GATE M9:GATE 823.354 
CC38394 M1:GATE M2:DRN 8.65e-18
CC38329 M1:GATE ZN:2 4.25e-18
CC38310 M1:GATE ZN:1 1.751e-17
CC38363 M9:GATE M10:DRN 4.597e-17
CC38309 M9:GATE ZN:1 8.55e-18
R15 M14:GATE I:5 111.3 
R16 M6:GATE I:5 86.5669 
R17 I I:5 23.5361 
R18 I:3 I:5 2065.9 
R19 I:4 I:5 21.0655 
R20 M13:GATE I:5 278.849 
R21 I:5 M5:GATE 235.694 
CC38382 I:5 M6:DRN 6.164e-17
CC38352 I:5 M14:DRN 1.64e-18
R22 M5:GATE M13:GATE 1058.4 
CC38377 M5:GATE M6:DRN 1.374e-17
CC38325 M5:GATE ZN:2 1.359e-17
CC38373 M13:GATE M6:DRN 1.28e-18
CC38347 M13:GATE M14:DRN 4.517e-17
CC38318 M13:GATE ZN:2 3.58e-18
CC38305 M13:GATE ZN:1 1.791e-17
R23 M15:GATE I:4 111.3 
R24 I I:4 23.2649 
R25 I:3 I:4 22.2029 
R26 I:4 M7:GATE 83.8364 
CC38371 I:4 M8:DRN 4.082e-17
CC38343 I:4 M16:DRN 1.58e-18
CC38367 M7:GATE M8:DRN 8.41e-18
CC38323 M7:GATE ZN:2 1.354e-17
R27 M8:GATE I:3 80.5597 
R28 I I:3 22.7377 
R29 I:3 M16:GATE 111.3 
CC38380 I:3 M6:DRN 1.555e-17
CC38370 I:3 M8:DRN 4.392e-17
CC38364 I:3 M10:DRN 1.306e-17
CC38395 I:3 M2:DRN 1.509e-17
CC38389 I:3 M4:DRN 1.533e-17
CC38331 I:3 ZN:2 5.526e-17
CC38358 I:3 M12:DRN 1.319e-17
CC38350 I:3 M14:DRN 1.335e-17
CC38342 I:3 M16:DRN 1.359e-17
CC38312 I:3 ZN:1 2.024e-17
CC38338 M16:GATE M16:DRN 4.714e-17
CC38302 M16:GATE ZN:1 6.15e-18
CC38379 I M6:DRN 1.45e-18
CC38369 I M8:DRN 2.28e-18
CC38330 I ZN:2 6.058e-17
CC38341 I M16:DRN 1.49e-18
CC38311 I ZN:1 5.424e-17
CC38386 M4:GATE M4:DRN 8.54e-18
CC38326 M4:GATE ZN:2 1.214e-17
CC38376 M6:GATE M6:DRN 8.54e-18
CC38324 M6:GATE ZN:2 1.42e-17
CC38366 M8:GATE M8:DRN 2.158e-17
CC38322 M8:GATE ZN:2 3.62e-18
CC38321 M10:GATE ZN:2 1.02e-18
CC38362 M10:GATE M10:DRN 4.502e-17
CC38308 M10:GATE ZN:1 1.839e-17
R30 M11:GATE M3:GATE 1074.97 
CC38320 M11:GATE ZN:2 7.92e-18
CC38356 M11:GATE M12:DRN 4.476e-17
CC38307 M11:GATE ZN:1 1.784e-17
CC38387 M3:GATE M4:DRN 1.204e-17
CC38327 M3:GATE ZN:2 1.501e-17
CC38355 M12:GATE M12:DRN 4.457e-17
CC38319 M12:GATE ZN:2 5.02e-18
CC38306 M12:GATE ZN:1 1.849e-17
CC38346 M14:GATE M14:DRN 4.563e-17
CC38304 M14:GATE ZN:1 1.787e-17
CC38339 M15:GATE M16:DRN 4.487e-17
CC38303 M15:GATE ZN:1 1.862e-17
CC38393 M2:GATE M2:DRN 8.41e-18
CC38328 M2:GATE ZN:2 8.1e-18
C31 I:1 0 5.64e-18
C32 I:2 0 6.533e-17
C33 M1:GATE 0 5.024e-17
C34 M9:GATE 0 1.0173e-16
C35 I:5 0 7.17e-18
C36 M5:GATE 0 3.067e-17
C37 M13:GATE 0 4.379e-17
C38 I:4 0 8.85e-18
C39 M7:GATE 0 3.415e-17
C40 I:3 0 1.091e-16
C41 M16:GATE 0 6.436e-17
C42 I 0 8.49e-17
C43 M4:GATE 0 3.199e-17
C44 M6:GATE 0 3.241e-17
C45 M8:GATE 0 2.877e-17
C46 M10:GATE 0 5.205e-17
C47 M11:GATE 0 4.88e-17
C48 M3:GATE 0 3.624e-17
C49 M12:GATE 0 4.186e-17
C50 M14:GATE 0 4.464e-17
C51 M15:GATE 0 5.667e-17
C52 M2:GATE 0 4.137e-17
R53 ZN:1 M12:DRN 14.9999 
R54 M12:DRN M11:SRC 0.001 
R55 M6:DRN ZN:2 15.181 
R56 M4:DRN ZN:2 14.9999 
R57 M8:DRN ZN:2 15.3164 
R58 ZN ZN:2 0.11093 
R59 ZN:2 M2:DRN 15.1433 
R60 M2:DRN M1:SRC 0.001 
R61 ZN ZN:1 0.09013 
R62 M16:DRN ZN:1 15.4792 
R63 M10:DRN ZN:1 15.1923 
R64 ZN:1 M14:DRN 15.3033 
R65 M16:DRN M14:DRN 1522.23 
R66 M14:DRN M13:SRC 0.001 
R67 M8:DRN M7:SRC 0.001 
R68 M10:DRN M9:SRC 0.001 
R69 M4:DRN M3:SRC 0.001 
R70 M6:DRN M5:SRC 0.001 
R71 M16:DRN M15:SRC 0.001 
C72 M12:DRN 0 3.99e-18
C73 ZN:2 0 1.788e-16
C74 M2:DRN 0 8.07e-18
C75 ZN 0 6.6e-19
C76 ZN:1 0 2.1896e-16
C77 M14:DRN 0 4e-18
C78 M8:DRN 0 8.97e-18
C79 M10:DRN 0 6.92e-18
C80 M4:DRN 0 5.42e-18
C81 M6:DRN 0 5.42e-18
C82 M16:DRN 0 6.06e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
