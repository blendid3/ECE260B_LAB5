.SUBCKT MUX2D1 I0 I1 S Z
MMM10 M7:DRN M10:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=7e-14  AS=5.3e-14  PD=9.55e-07  PS=7.25e-07  SA=3.08e-07  SB=4.3e-07  NRD=0.338  NRS=1.092  SCA=8.401  SCB=0.009  SCC=0.0006042 
MMM11 M7:SRC M11:GATE M8:DRN vdd pch L=6e-08 W=4.14e-07  AD=4.5e-14  AS=5.8e-14  PD=7.76e-07  PS=8.43e-07  SA=2.81e-07  SB=2.88e-07  NRD=1.953  NRS=0.397  SCA=6.236  SCB=0.006  SCC=0.0002084 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.9e-07  AD=6.8e-14  AS=5.1e-14  PD=1.13e-06  PS=6.5e-07  SA=6.31e-07  SB=1.75e-07  NRD=0.496  NRS=0.381  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=2.66e-07  AD=4.3e-14  AS=4.9e-14  PD=8.5e-07  PS=6.89e-07  SA=1.65e-07  SB=2.83e-07  NRD=0.72  NRS=0.87  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=5.1e-14  AS=4.2e-14  PD=6.5e-07  PS=7.3e-07  SA=2.52e-07  SB=4.95e-07  NRD=0.381  NRS=8.076  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=2.63e-07  AD=3.8e-14  AS=2.7e-14  PD=6.97e-07  PS=4.88e-07  SA=4.76e-07  SB=2.22e-07  NRD=0.581  NRS=7.566  SCA=15.388  SCB=0.017  SCC=0.002 
MMM4 M2:SRC M4:GATE M3:DRN vss nch L=6e-08 W=2.51e-07  AD=2.6e-14  AS=3.5e-14  PD=4.5e-07  PS=6.43e-07  SA=1.73e-07  SB=7.55e-07  NRD=0.473  NRS=0.622  SCA=5.308  SCB=0.005  SCC=6.294e-05 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=1.99e-07  AD=3.5e-14  AS=2e-14  PD=7.5e-07  PS=3.95e-07  SA=1.8e-07  SB=8.41e-07  NRD=0.972  NRS=0.553  SCA=13.679  SCB=0.016  SCC=0.001 
MMM6 vss M6:GATE M3:SRC vss nch L=6e-08 W=2.34e-07  AD=2.4e-14  AS=2.4e-14  PD=4.65e-07  PS=4.32e-07  SA=3.47e-07  SB=5.3e-07  NRD=9.028  NRS=1.899  SCA=13.049  SCB=0.015  SCC=0.001 
MMM7 M7:DRN M7:GATE M7:SRC vdd pch L=6e-08 W=3.43e-07  AD=4.6e-14  AS=3.8e-14  PD=6.25e-07  PS=6.44e-07  SA=3.36e-07  SB=7.6e-07  NRD=0.425  NRS=0.369  SCA=12.054  SCB=0.013  SCC=0.001 
MMM8 M8:DRN M8:GATE vdd vdd pch L=6e-08 W=3.17e-07  AD=4.4e-14  AS=5.8e-14  PD=6.37e-07  PS=8.21e-07  SA=2.54e-07  SB=4.6e-07  NRD=0.482  NRS=0.807  SCA=13.7  SCB=0.015  SCC=0.001 
MMM9 M9:DRN M9:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=8.6e-14  AS=5.3e-14  PD=1.37e-06  PS=7.25e-07  SA=6.86e-07  SB=1.65e-07  NRD=0.433  NRS=1.092  SCA=8.401  SCB=0.009  SCC=0.0006042 
R0 I0 M8:GATE 120.779 
R1 M8:GATE M6:GATE 361.546 
CC2981 M8:GATE M11:GATE 3.38e-18
CC2909 M8:GATE M12:DRN 6.6e-18
CC2996 M8:GATE S 1.342e-17
CC2989 M8:GATE M12:GATE 2.7e-18
CC2902 M8:GATE M8:DRN 3.652e-17
R2 M6:GATE I0 107.803 
CC2921 M6:GATE M3:GATE 1.87e-18
CC2915 M6:GATE M7:GATE 2.51e-18
CC2905 M6:GATE M3:SRC 1.038e-17
CC3007 M6:GATE M5:GATE 5.06e-18
CC2903 M6:GATE M8:DRN 3.84e-18
CC2923 I0 M3:GATE 1.51e-18
CC2917 I0 M7:GATE 4.52e-18
CC2911 I0 M12:DRN 1.568e-17
CC2906 I0 M3:SRC 8.642e-17
CC3013 I0 M5:GATE 4.15e-18
CC3001 I0 S 5.384e-17
CC2993 I0 M12:GATE 3.41e-18
CC2904 I0 M8:DRN 5.42e-18
C3 M8:GATE 0 3.584e-17
C4 M6:GATE 0 5.354e-17
C5 I0 0 1.462e-17
R6 M1:DRN Z 15.2788 
CC2929 M1:DRN M9:GATE 1.22e-18
CC2941 M1:DRN M1:GATE 2.197e-17
CC2950 M1:DRN M3:DRN 3.205e-17
R7 Z M9:DRN 15.4424 
CC2930 Z M9:GATE 1.579e-17
CC2972 Z I1 1.386e-17
CC2942 Z M1:GATE 1.145e-17
CC2951 Z M3:DRN 6.425e-17
CC2927 M9:DRN M9:GATE 4.818e-17
CC2934 M9:DRN M7:SRC 7.58e-18
C8 M1:DRN 0 2.617e-17
C9 Z 0 1.1794e-16
C10 M9:DRN 0 3.794e-17
R11 M1:GATE M9:GATE 421.02 
R12 M7:SRC M9:GATE 362.379 
R13 M9:GATE M3:DRN 375.433 
CC2963 M9:GATE I1 6.42e-18
CC2955 M9:GATE M10:GATE 5.76e-18
R14 M1:GATE M3:DRN 331.14 
R15 M3:DRN M7:SRC 74.1855 
CC3022 M3:DRN M4:GATE 2.35e-18
CC3019 M3:DRN M4:GATE 1.933e-17
CC3009 M3:DRN M5:GATE 8.3e-18
CC2966 M3:DRN I1 3.826e-17
CC2939 M3:DRN M7:GATE 1.7e-18
CC2946 M3:DRN M7:GATE 9.87e-18
CC2945 M3:DRN M7:DRN 1.97e-18
CC2944 M3:DRN M8:DRN 2.08e-18
CC2943 M3:DRN M12:DRN 1.868e-17
CC2948 M3:DRN M2:SRC 6.98e-17
CC2949 M3:DRN M3:GATE 3.276e-17
R16 M7:SRC M1:GATE 319.626 
CC3014 M7:SRC M4:GATE 3.53e-18
CC2953 M7:SRC M10:GATE 1.579e-17
CC2979 M7:SRC M11:GATE 3.74e-17
CC3004 M7:SRC M5:GATE 1.41e-18
CC2975 M7:SRC M2:GATE 1.01e-18
CC2938 M7:SRC M3:GATE 2.525e-17
CC2936 M7:SRC M3:SRC 5.645e-17
CC2935 M7:SRC M7:GATE 2.136e-17
CC2933 M7:SRC M7:DRN 5.138e-17
CC2932 M7:SRC M8:DRN 3.432e-17
CC2931 M7:SRC M12:DRN 1.972e-17
CC2959 M1:GATE M10:GATE 4.05e-18
CC2973 M1:GATE M2:GATE 1e-18
CC2970 M1:GATE I1 6.04e-18
CC2940 M1:GATE M12:DRN 4.268e-17
C17 M9:GATE 0 1.0921e-16
C18 M3:DRN 0 1.16e-17
C19 M7:SRC 0 3.707e-17
C20 M1:GATE 0 4.609e-17
R21 M7:DRN M2:SRC 60.9229 
CC2908 M7:DRN M12:DRN 7.41e-18
CC2913 M7:DRN M7:GATE 1.943e-17
CC2919 M7:DRN M3:GATE 1.528e-17
CC3015 M7:DRN M4:GATE 7.19e-18
CC2962 M7:DRN I1 6.266e-17
CC2954 M7:DRN M10:GATE 1.512e-17
CC2974 M7:DRN M2:GATE 3.62e-18
CC2916 M2:SRC M7:GATE 1.07e-18
CC2958 M2:SRC M10:GATE 2.56e-18
CC3020 M2:SRC M4:GATE 3.462e-17
CC2967 M2:SRC I1 3.23e-17
CC2976 M2:SRC M2:GATE 3.79e-18
C22 M7:DRN 0 8.21e-18
C23 M2:SRC 0 4.288e-17
R24 M2:GATE M10:GATE 585.413 
R25 M10:GATE I1 156.775 
CC2957 M10:GATE M7:GATE 5.49e-18
CC2952 M10:GATE M12:DRN 2.18e-18
R26 I1 M2:GATE 121.151 
CC2968 I1 M3:GATE 8e-18
C27 M10:GATE 0 7.907e-17
C28 I1 0 3.668e-17
C29 M2:GATE 0 6.292e-17
R30 M11:GATE M12:GATE 307.4 
R31 M5:GATE M12:GATE 604.588 
R32 M12:GATE S 190.285 
CC2985 M12:GATE M12:DRN 3.385e-17
CC2986 M12:GATE M8:DRN 6.13e-18
R33 S M5:GATE 104.362 
CC2999 S M5:DRN 7.595e-17
CC2994 S M12:DRN 2.07e-18
CC2995 S M8:DRN 2.88e-18
R34 M5:GATE M4:GATE 378.418 
CC3002 M5:GATE M12:DRN 1.551e-17
CC3003 M5:GATE M8:DRN 1.39e-18
CC3006 M5:GATE M3:SRC 5.11e-18
CC3008 M5:GATE M5:DRN 2.361e-17
CC3011 M5:GATE M3:GATE 3.54e-18
CC3021 M4:GATE M3:GATE 1.34e-18
CC3016 M4:GATE M7:GATE 3.27e-18
CC2977 M11:GATE M12:DRN 9.05e-18
CC2978 M11:GATE M8:DRN 2.578e-17
CC2982 M11:GATE M7:GATE 7.14e-18
C35 M12:GATE 0 1.2851e-16
C36 S 0 5.035e-17
C37 M5:GATE 0 1.3893e-16
C38 M4:GATE 0 6.027e-17
C39 M11:GATE 0 3.261e-17
R40 M8:DRN M3:SRC 60.9906 
CC2912 M8:DRN M7:GATE 1.143e-17
CC2907 M8:DRN M12:DRN 3.55e-17
CC2918 M8:DRN M3:GATE 2.87e-18
CC2920 M3:SRC M3:GATE 2.957e-17
C41 M8:DRN 0 2.551e-17
C42 M3:SRC 0 5.05e-18
R43 M12:DRN M7:GATE 203.264 
R44 M5:DRN M7:GATE 210.746 
R45 M7:GATE M3:GATE 250.426 
R46 M5:DRN M12:DRN 71.6841 
C47 M7:GATE 0 9.353e-17
C48 M3:GATE 0 6.4e-18
C49 M5:DRN 0 1.3972e-16
C50 M12:DRN 0 4.079e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
