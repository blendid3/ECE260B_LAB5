.SUBCKT XNR2D2 A1 A2 ZN
MMM10 M9:SRC M10:GATE vdd vdd pch L=6e-08 W=2.66e-07  AD=3.6e-14  AS=4.5e-14  PD=6.25e-07  PS=7.45e-07  SA=1.7e-07  SB=3.22e-07  NRD=0.561  NRS=0.684  SCA=15.255  SCB=0.017  SCC=0.002 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=2.64e-07  AD=4.5e-14  AS=4.2e-14  PD=7.45e-07  PS=8.4e-07  SA=1.6e-07  SB=1.75e-07  NRD=0.684  NRS=0.704  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7.2e-14  AS=3.9e-14  PD=1.15e-06  PS=5.9e-07  SA=8.63e-07  SB=1.85e-07  NRD=0.609  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 vdd M12:GATE M12:SRC vdd pch L=6e-08 W=5.24e-07  AD=7.8e-14  AS=5.2e-14  PD=1.34e-06  PS=7.2e-07  SA=1e-06  SB=1.5e-07  NRD=1.688  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=4.9e-14  PD=5.9e-07  PS=6.4e-07  SA=5.87e-07  SB=4.45e-07  NRD=4.141  NRS=0.654  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 M13:DRN M13:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.5e-14  PD=7.2e-07  PS=7.7e-07  SA=7.09e-07  SB=4.1e-07  NRD=2.099  NRS=0.66  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=4.9e-14  AS=4.2e-14  PD=6.4e-07  PS=7.48e-07  SA=2.3e-07  SB=7.55e-07  NRD=0.654  NRS=8.791  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M8:SRC M14:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.7e-14  AS=6.5e-14  PD=8.53e-07  PS=7.7e-07  SA=3.1e-07  SB=7.2e-07  NRD=4.762  NRS=0.66  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE M4:SRC vss nch L=6e-08 W=1.95e-07  AD=3e-14  AS=1.9e-14  PD=5.63e-07  PS=3.9e-07  SA=6.26e-07  SB=1.99e-07  NRD=0.843  NRS=8.478  SCA=18.359  SCB=0.02  SCC=0.002 
MMM5 M3:SRC M5:GATE M4:DRN vss nch L=6e-08 W=2.36e-07  AD=2.4e-14  AS=3.6e-14  PD=4.32e-07  PS=6.67e-07  SA=1.74e-07  SB=1.015e-06  NRD=0.499  NRS=0.721  SCA=6.258  SCB=0.006  SCC=0.0001231 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=1.99e-07  AD=3.4e-14  AS=2.2e-14  PD=7.4e-07  PS=4.46e-07  SA=1.75e-07  SB=4.11e-07  NRD=0.947  NRS=1.704  SCA=13.679  SCB=0.016  SCC=0.001 
MMM7 M4:SRC M7:GATE vss vss nch L=6.2e-08 W=1.92e-07  AD=1.9e-14  AS=2.1e-14  PD=3.9e-07  PS=4.34e-07  SA=3.39e-07  SB=4.78e-07  NRD=8.478  NRS=0.609  SCA=18.359  SCB=0.02  SCC=0.002 
MMM8 M8:DRN M8:GATE M8:SRC vdd pch L=6e-08 W=3.72e-07  AD=3.9e-14  AS=4e-14  PD=6.97e-07  PS=6.07e-07  SA=2.64e-07  SB=9.9e-07  NRD=10.154  NRS=0.34  SCA=12.196  SCB=0.013  SCC=0.001 
MMM9 M8:DRN M9:GATE M9:SRC vdd pch L=6e-08 W=2.4e-07  AD=2.5e-14  AS=3.3e-14  PD=4.43e-07  PS=5.65e-07  SA=2.46e-07  SB=1.25e-06  NRD=0.476  NRS=0.612  SCA=6.833  SCB=0.007  SCC=0.000198 
R0 M4:SRC M9:SRC 60.6379 
CC29572 M4:SRC M6:GATE 2.84e-18
CC29617 M4:SRC M8:DRN 7.123e-17
CC29513 M4:SRC M4:GATE 3.081e-17
CC29521 M4:SRC M10:GATE 2.043e-17
CC29524 M4:SRC M7:GATE 1.004e-17
CC29529 M4:SRC M3:SRC 3.043e-17
CC29586 M9:SRC N_12:1 1.68e-18
CC29634 M9:SRC M4:DRN 1.9e-18
CC29551 M9:SRC M11:GATE 3.46e-18
CC29510 M9:SRC M8:GATE 8.33e-18
CC29508 M9:SRC M11:SRC 4.178e-17
CC29512 M9:SRC M4:GATE 2.01e-18
CC29519 M9:SRC M10:GATE 3.996e-17
CC29522 M9:SRC M7:GATE 4.88e-18
CC29562 M9:SRC A1 2.255e-17
CC29557 M9:SRC M9:GATE 2.36e-17
C1 M4:SRC 0 6.44e-18
C2 M9:SRC 0 1.605e-17
R3 M5:GATE M6:GATE 383.19 
CC29640 M5:GATE M4:DRN 2.641e-17
CC29576 M5:GATE M8:GATE 3.35e-18
CC29618 M5:GATE M8:DRN 2.12e-18
CC29579 M5:GATE M3:SRC 4.606e-17
CC29580 M5:GATE M4:GATE 1.63e-18
R4 A1 M6:GATE 96.8281 
R5 M6:GATE M11:GATE 583.368 
CC29568 M6:GATE M11:SRC 1.602e-17
CC29575 M6:GATE M4:GATE 2.87e-18
CC29574 M6:GATE M3:SRC 1.967e-17
CC29573 M6:GATE M6:DRN 3.108e-17
R6 M9:GATE M11:GATE 317.206 
R7 M11:GATE A1 199.983 
CC29549 M11:GATE M11:SRC 2.931e-17
CC29550 M11:GATE M10:GATE 1.04e-18
CC29584 M11:GATE N_12:1 2.18e-18
CC29564 A1 M7:GATE 1.509e-17
CC29566 A1 M6:DRN 6.785e-17
CC29560 A1 M11:SRC 7.67e-18
CC29561 A1 M10:GATE 5.24e-18
CC29555 M9:GATE M11:SRC 1.466e-17
CC29556 M9:GATE M10:GATE 3.2e-18
CC29558 M9:GATE M8:GATE 5.95e-18
CC29615 M9:GATE M8:DRN 3.408e-17
CC29587 M9:GATE N_12:1 2.69e-18
C8 M5:GATE 0 5.181e-17
C9 M6:GATE 0 1.3845e-16
C10 M11:GATE 0 1.2697e-16
C11 A1 0 7.396e-17
C12 M9:GATE 0 3.276e-17
R13 M4:GATE M8:GATE 230.551 
CC29642 M4:GATE M4:DRN 2.504e-17
CC29620 M4:GATE M8:DRN 2.861e-17
CC29517 M4:GATE M8:SRC 9.58e-18
CC29536 M4:GATE M14:GATE 2.33e-18
CC29530 M4:GATE M3:SRC 1.337e-17
CC29548 M4:GATE M3:GATE 4.96e-18
R14 M6:DRN M8:GATE 218.1 
R15 M8:GATE M11:SRC 211.21 
CC29588 M8:GATE N_12:1 1.991e-17
CC29636 M8:GATE M4:DRN 2.292e-17
CC29616 M8:GATE M8:DRN 1.9e-18
CC29523 M8:GATE M7:GATE 4.28e-18
CC29516 M8:GATE M8:SRC 2.347e-17
CC29534 M8:GATE M14:GATE 3.23e-18
CC29528 M8:GATE M3:SRC 2.28e-18
R16 M11:SRC M6:DRN 71.0738 
CC29632 M11:SRC M4:DRN 4.879e-17
CC29611 M11:SRC M8:DRN 1.392e-17
CC29518 M11:SRC M10:GATE 5.23e-18
CC29514 M11:SRC M8:SRC 5.64e-18
CC29533 M11:SRC M14:GATE 2.66e-18
CC29527 M11:SRC M3:SRC 1.82e-18
C17 M4:GATE 0 1.134e-17
C18 M8:GATE 0 8.823e-17
C19 M11:SRC 0 5.469e-17
C20 M6:DRN 0 1.3609e-16
R21 M1:SRC M2:DRN 0.001 
R22 M2:DRN ZN 15.4947 
CC29595 M2:DRN N_12:1 8.732e-17
CC29543 M2:DRN A2 1.11e-18
CC29625 M2:DRN M1:GATE 1.046e-17
CC29629 M2:DRN M2:GATE 1.189e-17
R23 ZN M12:SRC 30.6142 
CC29643 ZN M4:DRN 5.563e-17
CC29603 ZN M13:GATE 3.56e-18
CC29624 ZN M1:GATE 1.334e-17
CC29627 ZN M2:GATE 3.84e-18
CC29607 ZN M12:GATE 2.784e-17
CC29544 ZN A2 1.42e-17
CC29596 ZN N_12:1 1.274e-17
R24 M12:SRC M13:DRN 0.001 
CC29583 M12:SRC N_12:1 6.37e-18
CC29606 M12:SRC M12:GATE 3.134e-17
CC29600 M12:SRC M13:GATE 2.804e-17
C25 M2:DRN 0 1.066e-17
C26 ZN 0 1.2423e-16
C27 M12:SRC 0 5.89e-18
R28 M10:GATE M7:GATE 139.125 
R29 M3:SRC M7:GATE 162.608 
R30 M7:GATE M8:SRC 167.452 
CC29589 M7:GATE N_12:1 4.411e-17
CC29637 M7:GATE M4:DRN 1.4e-18
R31 M8:SRC M3:SRC 74.6692 
CC29582 M8:SRC N_12:1 7.545e-17
CC29531 M8:SRC M14:GATE 1.94e-17
CC29539 M8:SRC A2 1.185e-17
CC29542 M3:SRC A2 7.063e-17
CC29641 M3:SRC M4:DRN 6.33e-18
CC29619 M3:SRC M8:DRN 5.05e-18
CC29547 M3:SRC M3:GATE 1.501e-17
CC29535 M3:SRC M14:GATE 5.87e-18
C32 M10:GATE 0 3.437e-17
C33 M7:GATE 0 6.686e-17
C34 M8:SRC 0 8.174e-17
C35 M3:SRC 0 8.99e-18
R36 A2 M14:GATE 152.373 
R37 M14:GATE M3:GATE 545.918 
CC29581 M14:GATE N_12:1 1.752e-17
CC29598 M14:GATE M13:GATE 4.54e-18
R38 M3:GATE A2 118.665 
CC29594 M3:GATE N_12:1 4.46e-18
CC29597 A2 N_12:1 2.46e-18
CC29604 A2 M13:GATE 1.04e-18
CC29608 A2 M12:GATE 2.33e-18
CC29622 A2 M8:DRN 3.891e-17
CC29626 A2 M2:GATE 2.59e-18
CC29644 A2 M4:DRN 2.13e-18
C39 M14:GATE 0 7.238e-17
C40 M3:GATE 0 5.095e-17
C41 A2 0 4.936e-17
R42 N_12:1 M12:GATE 149.883 
R43 M12:GATE M1:GATE 680.901 
R44 M1:GATE N_12:1 144.19 
R45 M13:GATE N_12:1 104.675 
R46 M4:DRN N_12:1 79.1803 
R47 M8:DRN N_12:1 76.881 
R48 N_12:1 M2:GATE 88.5713 
R49 M8:DRN M4:DRN 99.8668 
C50 M12:GATE 0 5.266e-17
C51 M1:GATE 0 5.75e-17
C52 N_12:1 0 3.534e-17
C53 M2:GATE 0 4.677e-17
C54 M8:DRN 0 1.457e-17
C55 M4:DRN 0 2.678e-17
C56 M13:GATE 0 5.75e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
