.SUBCKT INVD24 I ZN
MMM20 M20:DRN M20:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.2e-06  SB=5e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM21 vss M21:GATE M21:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.4e-07  SB=5.26e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM22 M22:DRN M22:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=5.52e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM23 vss M23:GATE M23:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=5.78e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM24 vss M24:GATE M24:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.6e-07  SB=6.04e-06  NRD=0.567  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM25 vdd M25:GATE M25:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=6.04e-06  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM26 M26:DRN M26:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=5.78e-06  SB=4.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM27 vdd M27:GATE M27:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=5.54e-06  SB=6.6e-07  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM28 M28:DRN M28:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=5.28e-06  SB=9.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM29 vdd M29:GATE M29:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=5.04e-06  SB=1.16e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM40 M40:DRN M40:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.24e-06  SB=3.96e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM41 vdd M41:GATE M41:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.98e-06  SB=4.22e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM42 M42:DRN M42:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.72e-06  SB=4.48e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM43 vdd M43:GATE M43:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.46e-06  SB=4.74e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM44 M44:DRN M44:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.2e-06  SB=5e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM45 vdd M45:GATE M45:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.4e-07  SB=5.26e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM46 M46:DRN M46:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=5.52e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM47 vdd M47:GATE M47:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=5.78e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=3.78e-06  SB=2.42e-06  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM48 M48:DRN M48:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=6.04e-06  NRD=2.057  NRS=0.532  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=3.54e-06  SB=2.66e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=6.04e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.28e-06  SB=2.92e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=5.78e-06  SB=4.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=3.02e-06  SB=3.18e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=5.54e-06  SB=6.6e-07  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.76e-06  SB=3.44e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=5.28e-06  SB=9.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vss M15:GATE M15:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.5e-06  SB=3.7e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=5.04e-06  SB=1.16e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.24e-06  SB=3.96e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=4.78e-06  SB=1.42e-06  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 vss M17:GATE M17:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.98e-06  SB=4.22e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=4.54e-06  SB=1.66e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M18:DRN M18:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.72e-06  SB=4.48e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=4.28e-06  SB=1.92e-06  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vss M19:GATE M19:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.46e-06  SB=4.74e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=4.04e-06  SB=2.16e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM30 M30:DRN M30:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=4.78e-06  SB=1.42e-06  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM31 vdd M31:GATE M31:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=4.54e-06  SB=1.66e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM32 M32:DRN M32:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=4.28e-06  SB=1.92e-06  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM33 vdd M33:GATE M33:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=4.04e-06  SB=2.16e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM34 M34:DRN M34:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=3.78e-06  SB=2.42e-06  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM35 vdd M35:GATE M35:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=3.54e-06  SB=2.66e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM36 M36:DRN M36:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=3.25e-06  SB=2.91e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM37 vdd M37:GATE M37:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.99e-06  SB=3.17e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM38 M38:DRN M38:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.76e-06  SB=3.44e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM39 vdd M39:GATE M39:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.5e-06  SB=3.7e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 I:24 I:6 22.6864 
R1 I:18 I:6 42.2554 
R2 I:7 I:6 0.69233 
R3 I:12 I:6 26.8311 
R4 I:6 I:17 17.5848 
CC15492 I:6 ZN:6 2.1131e-16
CC15540 I:6 ZN:7 1.624e-16
CC15414 I:6 ZN:1 1.383e-17
CC15666 I:6 M40:DRN 1.61e-18
CC15719 I:6 M22:DRN 1.39e-18
CC15740 I:6 M18:DRN 1.39e-18
CC15730 I:6 M20:DRN 1.39e-18
CC15690 I:6 M42:DRN 1.61e-18
CC15684 I:6 M44:DRN 1.61e-18
CC15678 I:6 M46:DRN 1.61e-18
CC15672 I:6 M48:DRN 1.58e-18
CC15708 I:6 M24:SRC 1.15e-18
CC15698 I:6 M16:DRN 1.39e-18
R5 M16:GATE I:17 81.2035 
R6 M40:GATE I:17 98.4282 
R7 I:24 I:17 22.2191 
R8 I:17 I:12 36.2001 
CC15493 I:17 ZN:6 2.05e-18
CC15699 I:17 M16:DRN 4.077e-17
R9 M41:GATE I:12 111.3 
R10 M17:GATE I:12 94.0755 
R11 I:18 I:12 37.0531 
R12 I:12 I:7 139.907 
CC15491 I:12 ZN:6 1.12e-18
CC15739 I:12 M18:DRN 3.736e-17
R13 I:25 I:7 22 
R14 I:18 I:7 29.085 
R15 I:26 I:7 33.2849 
R16 I:8 I:7 0.69344 
R17 I:7 I:27 66.914 
R18 M21:GATE I:27 82.8124 
R19 M45:GATE I:27 100.037 
R20 I:13 I:27 34.0521 
R21 I:26 I:27 21.9048 
R22 I:27 I:8 24.5967 
CC15717 I:27 M22:DRN 4.061e-17
R23 I:14 I:8 108.561 
R24 I:9 I:8 0.45783 
R25 I:13 I:8 29.306 
R26 I:8 I:26 66.914 
R27 M44:GATE I:26 103.792 
R28 I:25 I:26 21.5119 
R29 I:26 M20:GATE 86.5669 
CC15488 I:26 ZN:6 1.26e-18
CC15727 I:26 M20:DRN 4.077e-17
CC15463 M20:GATE ZN:6 1.566e-17
CC15721 M20:GATE M20:DRN 4.57e-18
R30 M18:GATE I:18 80.5597 
R31 M42:GATE I:18 97.7846 
R32 I:18 I:25 22.4472 
CC15490 I:18 ZN:6 1.26e-18
CC15738 I:18 M18:DRN 4.077e-17
R33 M43:GATE I:25 101.061 
R34 I:25 M19:GATE 83.8364 
CC15728 I:25 M20:DRN 4.067e-17
CC15464 M19:GATE ZN:6 1.406e-17
CC15722 M19:GATE M20:DRN 4.57e-18
R35 M22:GATE I:13 94.0755 
R36 M46:GATE I:13 111.3 
R37 I:14 I:13 30.993 
R38 I:13 I:9 117.247 
CC15486 I:13 ZN:6 1.32e-18
CC15716 I:13 M22:DRN 3.9e-17
R39 M24:GATE I:9 466.584 
R40 I I:9 0.3368 
R41 I:14 I:9 25.7917 
R42 I:9 M48:GATE 552.017 
CC15705 I:9 M24:SRC 8.4e-18
R43 M24:GATE M48:GATE 686.528 
R44 M48:GATE I:14 222.947 
CC15506 M48:GATE ZN:7 5.1e-18
CC15458 M48:GATE ZN:6 4.04e-18
CC15667 M48:GATE M48:DRN 4.595e-17
R45 M24:GATE I:14 188.443 
R46 M47:GATE I:14 111.3 
R47 I:14 M23:GATE 94.0755 
CC15706 I:14 M24:SRC 3.854e-17
CC15460 M23:GATE ZN:6 1.376e-17
CC15701 M23:GATE M24:SRC 6.81e-18
R48 M39:GATE I:24 88.7752 
R49 M15:GATE I:24 94.0755 
R50 I:2 I:24 57.4715 
R51 M14:GATE I:24 222.334 
R52 I:24 M38:GATE 263.044 
CC15484 I:24 ZN:6 9.224e-17
CC15571 I:24 M34:DRN 1.114e-17
CC15565 I:24 M36:DRN 1.105e-17
CC15559 I:24 M38:DRN 1.097e-17
CC15589 I:24 M28:DRN 1.114e-17
CC15583 I:24 M30:DRN 1.114e-17
CC15577 I:24 M32:DRN 1.114e-17
CC15532 I:24 ZN:7 6.235e-17
CC15413 I:24 ZN:1 3.777e-17
CC15648 I:24 M4:DRN 1.643e-17
CC15638 I:24 M6:DRN 1.643e-17
CC15665 I:24 M40:DRN 1.114e-17
CC15657 I:24 M2:DRN 1.614e-17
CC15609 I:24 M12:DRN 1.632e-17
CC15601 I:24 M14:DRN 2.798e-17
CC15594 I:24 M26:DRN 1.097e-17
CC15628 I:24 M8:DRN 1.643e-17
CC15618 I:24 M10:DRN 1.643e-17
CC15725 I:24 M20:DRN 1.643e-17
CC15714 I:24 M22:DRN 1.643e-17
CC15736 I:24 M18:DRN 1.643e-17
CC15689 I:24 M42:DRN 1.114e-17
CC15683 I:24 M44:DRN 1.114e-17
CC15677 I:24 M46:DRN 1.114e-17
CC15671 I:24 M48:DRN 1.105e-17
CC15704 I:24 M24:SRC 1.614e-17
CC15696 I:24 M16:DRN 4.042e-17
R53 I:2 M38:GATE 284.964 
R54 M38:GATE M14:GATE 1102.4 
CC15556 M38:GATE M38:DRN 4.517e-17
CC15516 M38:GATE ZN:7 1.468e-17
CC15396 M38:GATE ZN:1 1.07e-18
CC15596 M38:GATE M14:DRN 3.25e-18
R55 M14:GATE I:2 240.862 
CC15469 M14:GATE ZN:6 1.279e-17
CC15598 M14:GATE M14:DRN 1.665e-17
R56 M37:GATE I:2 111.3 
R57 M36:GATE I:2 275.689 
R58 M12:GATE I:2 233.022 
R59 M13:GATE I:2 94.0755 
R60 I:2 I:3 60.2341 
CC15415 I:2 ZN:1 6.94e-18
CC15610 I:2 M12:DRN 1.33e-17
CC15603 I:2 M14:DRN 4.648e-17
R61 M35:GATE I:3 111.3 
R62 M36:GATE I:3 275.689 
R63 M12:GATE I:3 233.022 
R64 M11:GATE I:3 94.0755 
R65 I:16 I:3 31.8091 
R66 I:3 I:10 41.7693 
CC15495 I:3 ZN:6 1.41e-18
CC15611 I:3 M12:DRN 5.861e-17
R67 I:16 I:10 18.5804 
R68 I:20 I:10 22 
R69 I:21 I:10 44.2281 
R70 I:5 I:10 0.45838 
R71 I:10 I:19 22.6293 
CC15499 I:10 ZN:6 2.0845e-16
CC15590 I:10 M28:DRN 1.6e-18
CC15584 I:10 M30:DRN 1.6e-18
CC15578 I:10 M32:DRN 1.6e-18
CC15572 I:10 M34:DRN 1.6e-18
CC15546 I:10 ZN:7 1.6008e-16
CC15420 I:10 ZN:1 1.372e-17
CC15649 I:10 M4:DRN 1.31e-18
CC15639 I:10 M6:DRN 1.31e-18
CC15658 I:10 M2:DRN 1.07e-18
CC15595 I:10 M26:DRN 1.52e-18
CC15631 I:10 M8:DRN 1.31e-18
CC15623 I:10 M10:DRN 1.31e-18
R72 I:16 I:19 22.1694 
R73 M9:GATE I:19 85.0652 
R74 I:20 I:19 21.0442 
R75 I:19 M33:GATE 111.3 
CC15497 I:19 ZN:6 1.41e-18
CC15621 I:19 M10:DRN 4.003e-17
CC15569 M33:GATE M34:DRN 4.48e-17
CC15521 M33:GATE ZN:7 1.782e-17
CC15483 I ZN:6 4.4e-18
CC15531 I ZN:7 8.14e-18
R76 I:23 M1:GATE 133.769 
R77 M1:GATE M25:GATE 692.112 
CC15482 M1:GATE ZN:6 3.89e-18
CC15656 M1:GATE M2:DRN 8.28e-18
R78 M25:GATE I:23 158.262 
CC15529 M25:GATE ZN:7 4.91e-18
CC15593 M25:GATE M26:DRN 4.573e-17
R79 M26:GATE I:23 111.3 
R80 M2:GATE I:23 82.8124 
R81 I:15 I:23 21.3025 
R82 I:23 I:11 22.6864 
CC15505 I:23 ZN:6 2.73e-18
CC15660 I:23 M2:DRN 7.86e-17
R83 I:5 I:11 0.69092 
R84 I:1 I:11 51.3138 
R85 I:4 I:11 28.2443 
R86 I:11 I:15 17.5848 
R87 M27:GATE I:15 111.3 
R88 M3:GATE I:15 81.2035 
R89 I:15 I:4 36.2001 
CC15504 I:15 ZN:6 2.26e-18
CC15652 I:15 M4:DRN 4.143e-17
R90 M28:GATE I:4 111.3 
R91 M4:GATE I:4 94.0755 
R92 I:5 I:4 160.59 
R93 I:4 I:1 28.0967 
CC15503 I:4 ZN:6 1.43e-18
CC15651 I:4 M4:DRN 3.759e-17
R94 M29:GATE I:1 111.3 
R95 M5:GATE I:1 94.0755 
R96 I:22 I:1 35.1071 
R97 I:1 I:5 45.9733 
CC15502 I:1 ZN:6 1.41e-18
CC15642 I:1 M6:DRN 3.716e-17
R98 I:21 I:5 44.2281 
R99 I:5 I:22 17.575 
R100 M30:GATE I:22 111.3 
R101 I:21 I:22 21.5119 
R102 I:22 M6:GATE 81.9458 
CC15501 I:22 ZN:6 2.54e-18
CC15641 I:22 M6:DRN 4.03e-17
CC15477 M6:GATE ZN:6 1.179e-17
CC15635 M6:GATE M6:DRN 4.57e-18
CC15481 M2:GATE ZN:6 1.136e-17
CC15655 M2:GATE M2:DRN 4.59e-18
CC15480 M3:GATE ZN:6 1.204e-17
CC15646 M3:GATE M4:DRN 4.57e-18
CC15479 M4:GATE ZN:6 1.29e-17
CC15645 M4:GATE M4:DRN 7.44e-18
CC15478 M5:GATE ZN:6 1.29e-17
CC15636 M5:GATE M6:DRN 7.91e-18
R103 M7:GATE I:21 83.8364 
CC15476 M7:GATE ZN:6 1.29e-17
CC15626 M7:GATE M8:DRN 4.57e-18
R104 M31:GATE I:21 111.3 
R105 I:21 I:20 21.5119 
CC15500 I:21 ZN:6 1.41e-18
CC15632 I:21 M8:DRN 4.046e-17
R106 M8:GATE I:20 86.5669 
R107 I:20 M32:GATE 111.3 
CC15498 I:20 ZN:6 1.43e-18
CC15630 I:20 M8:DRN 4.011e-17
CC15574 M32:GATE M32:DRN 4.47e-17
CC15522 M32:GATE ZN:7 1.677e-17
CC15475 M8:GATE ZN:6 1.29e-17
CC15625 M8:GATE M8:DRN 5.62e-18
CC15474 M9:GATE ZN:6 1.29e-17
CC15616 M9:GATE M10:DRN 4.94e-18
CC15512 M42:GATE ZN:7 1.852e-17
CC15686 M42:GATE M42:DRN 4.557e-17
CC15511 M43:GATE ZN:7 1.669e-17
CC15681 M43:GATE M44:DRN 4.492e-17
CC15510 M44:GATE ZN:7 1.852e-17
CC15680 M44:GATE M44:DRN 4.557e-17
CC15509 M45:GATE ZN:7 1.669e-17
CC15675 M45:GATE M46:DRN 4.488e-17
CC15508 M46:GATE ZN:7 1.854e-17
CC15674 M46:GATE M46:DRN 4.557e-17
CC15507 M47:GATE ZN:7 1.649e-17
CC15668 M47:GATE M48:DRN 4.484e-17
R108 M10:GATE I:16 81.2035 
R109 I:16 M34:GATE 111.3 
CC15496 I:16 ZN:6 2.05e-18
CC15620 I:16 M10:DRN 4.117e-17
CC15568 M34:GATE M34:DRN 4.47e-17
CC15520 M34:GATE ZN:7 1.677e-17
CC15466 M17:GATE ZN:6 1.253e-17
CC15733 M17:GATE M18:DRN 8.21e-18
CC15700 M24:GATE M24:SRC 3.795e-17
CC15470 M13:GATE ZN:6 1.078e-17
CC15410 M13:GATE ZN:1 1.22e-18
CC15599 M13:GATE M14:DRN 1.36e-17
CC15514 M40:GATE ZN:7 1.713e-17
CC15662 M40:GATE M40:DRN 4.557e-17
CC15513 M41:GATE ZN:7 1.603e-17
CC15687 M41:GATE M42:DRN 4.516e-17
CC15473 M10:GATE ZN:6 1.228e-17
CC15615 M10:GATE M10:DRN 4.57e-18
CC15472 M11:GATE ZN:6 1.24e-17
CC15607 M11:GATE M12:DRN 5.62e-18
R110 M12:GATE M36:GATE 1066.52 
CC15471 M12:GATE ZN:6 1.166e-17
CC15411 M12:GATE ZN:1 3.76e-18
CC15606 M12:GATE M12:DRN 1.4e-17
CC15562 M36:GATE M36:DRN 4.495e-17
CC15518 M36:GATE ZN:7 1.556e-17
CC15398 M36:GATE ZN:1 4.98e-18
CC15468 M15:GATE ZN:6 2.2e-18
CC15693 M15:GATE M16:DRN 2.186e-17
CC15467 M16:GATE ZN:6 1.217e-17
CC15692 M16:GATE M16:DRN 4.57e-18
CC15465 M18:GATE ZN:6 1.566e-17
CC15732 M18:GATE M18:DRN 4.57e-18
CC15462 M21:GATE ZN:6 1.406e-17
CC15711 M21:GATE M22:DRN 4.57e-18
CC15461 M22:GATE ZN:6 1.563e-17
CC15710 M22:GATE M22:DRN 6.34e-18
CC15563 M35:GATE M36:DRN 4.475e-17
CC15519 M35:GATE ZN:7 1.782e-17
CC15557 M37:GATE M38:DRN 4.49e-17
CC15517 M37:GATE ZN:7 1.485e-17
CC15397 M37:GATE ZN:1 6.04e-18
CC15515 M39:GATE ZN:7 1.486e-17
CC15395 M39:GATE ZN:1 1.77e-18
CC15663 M39:GATE M40:DRN 4.547e-17
CC15587 M27:GATE M28:DRN 4.524e-17
CC15527 M27:GATE ZN:7 1.776e-17
CC15528 M26:GATE ZN:7 1.661e-17
CC15592 M26:GATE M26:DRN 4.461e-17
CC15586 M28:GATE M28:DRN 4.459e-17
CC15526 M28:GATE ZN:7 1.677e-17
CC15581 M29:GATE M30:DRN 4.468e-17
CC15525 M29:GATE ZN:7 1.782e-17
CC15580 M30:GATE M30:DRN 4.456e-17
CC15524 M30:GATE ZN:7 1.677e-17
CC15575 M31:GATE M32:DRN 4.48e-17
CC15523 M31:GATE ZN:7 1.782e-17
C111 I:6 0 1.129e-17
C112 I:17 0 7.39e-18
C113 I:12 0 2.6e-18
C114 I:7 0 8.35e-18
C115 I:27 0 4.56e-18
C116 I:8 0 1.052e-17
C117 I:26 0 3.86e-18
C118 M20:GATE 0 1.953e-17
C119 I:18 0 6.36e-18
C120 I:25 0 3.9e-18
C121 M19:GATE 0 2.316e-17
C122 I:13 0 2.84e-18
C123 I:9 0 8.48e-18
C124 M48:GATE 0 6.816e-17
C125 I:14 0 2.961e-17
C126 M23:GATE 0 3.215e-17
C127 I:24 0 2.0339e-16
C128 M38:GATE 0 2.66e-18
C129 M14:GATE 0 1.368e-17
C130 I:2 0 1.03e-18
C131 I:3 0 2.6e-18
C132 I:10 0 9.29e-18
C133 I:19 0 6.84e-18
C134 M33:GATE 0 2.83e-17
C135 I 0 6.27e-17
C136 M1:GATE 0 6.374e-17
C137 M25:GATE 0 8.776e-17
C138 I:23 0 1.018e-17
C139 I:11 0 1.668e-17
C140 I:15 0 2.38e-18
C141 I:4 0 2.79e-18
C142 I:1 0 2.85e-18
C143 I:5 0 1.053e-17
C144 I:22 0 2.81e-18
C145 M6:GATE 0 2.328e-17
C146 M2:GATE 0 3.259e-17
C147 M3:GATE 0 2.405e-17
C148 M4:GATE 0 2.895e-17
C149 M5:GATE 0 2.222e-17
C150 M7:GATE 0 2.28e-17
C151 I:21 0 2.92e-18
C152 I:20 0 2.81e-18
C153 M32:GATE 0 3.476e-17
C154 M8:GATE 0 2.838e-17
C155 M9:GATE 0 2.235e-17
C156 M42:GATE 0 3.939e-17
C157 M43:GATE 0 3.402e-17
C158 M44:GATE 0 3.238e-17
C159 M45:GATE 0 3.471e-17
C160 M46:GATE 0 4.121e-17
C161 M47:GATE 0 3.936e-17
C162 I:16 0 1.394e-17
C163 M34:GATE 0 2.881e-17
C164 M17:GATE 0 2.264e-17
C165 M24:GATE 0 2.792e-17
C166 M13:GATE 0 1.326e-17
C167 M40:GATE 0 3.418e-17
C168 M41:GATE 0 3.215e-17
C169 M10:GATE 0 2.239e-17
C170 M11:GATE 0 2.795e-17
C171 M12:GATE 0 2.019e-17
C172 M36:GATE 0 6.63e-18
C173 M15:GATE 0 2.557e-17
C174 M16:GATE 0 2.303e-17
C175 M18:GATE 0 2.523e-17
C176 M21:GATE 0 2.296e-17
C177 M22:GATE 0 2.946e-17
C178 M35:GATE 0 2.053e-17
C179 M37:GATE 0 3.29e-18
C180 M39:GATE 0 3.703e-17
C181 M27:GATE 0 3.055e-17
C182 M26:GATE 0 3.818e-17
C183 M28:GATE 0 3.491e-17
C184 M29:GATE 0 2.849e-17
C185 M30:GATE 0 2.907e-17
C186 M31:GATE 0 2.925e-17
R187 M21:SRC M22:DRN 0.001 
R188 ZN:5 M22:DRN 15.9319 
R189 M20:DRN M22:DRN 1282.24 
R190 M22:DRN M24:SRC 645.076 
R191 ZN:5 M24:SRC 16.1299 
R192 M20:DRN M24:SRC 1298.17 
R193 M24:SRC M23:SRC 0.001 
R194 ZN:3 M42:DRN 14.9999 
R195 M42:DRN M41:SRC 0.001 
R196 M31:SRC M32:DRN 0.001 
R197 M32:DRN ZN:2 14.9999 
R198 M34:DRN ZN:2 24.4354 
R199 M36:DRN ZN:2 63.8776 
R200 M28:DRN ZN:2 15.868 
R201 M30:DRN ZN:2 15.4503 
R202 M26:DRN ZN:2 16.0517 
R203 ZN:2 ZN:1 0.46131 
R204 ZN ZN:1 0.104 
R205 M38:DRN ZN:1 14.9999 
R206 M34:DRN ZN:1 39.8599 
R207 M36:DRN ZN:1 19.7443 
R208 ZN:3 ZN:1 0.436 
R209 ZN:1 M40:DRN 36.2236 
R210 ZN:3 M40:DRN 25.9096 
R211 M40:DRN M39:SRC 0.001 
R212 M48:DRN ZN:7 14.9999 
R213 M44:DRN ZN:7 45.7243 
R214 M46:DRN ZN:7 22.5904 
R215 ZN:7 ZN:3 0.55035 
R216 M44:DRN ZN:3 22.7254 
R217 ZN:3 M46:DRN 45.7243 
R218 M46:DRN M45:SRC 0.001 
R219 M25:SRC M26:DRN 0.001 
R220 M28:DRN M26:DRN 689.48 
R221 M26:DRN M30:DRN 835.354 
R222 M30:DRN M29:SRC 0.001 
R223 M28:DRN M27:SRC 0.001 
R224 M44:DRN M43:SRC 0.001 
R225 M48:DRN M47:SRC 0.001 
R226 ZN:5 M16:DRN 25.0067 
R227 ZN:6 M16:DRN 38.196 
R228 M16:DRN M15:SRC 0.001 
R229 M35:SRC M36:DRN 0.001 
R230 M13:SRC M14:DRN 0.001 
R231 M14:DRN ZN:6 14.9999 
R232 M12:DRN ZN:6 15.0192 
R233 M8:DRN ZN:6 47.6061 
R234 ZN:5 ZN:6 0.47459 
R235 ZN ZN:6 0.10123 
R236 M10:DRN ZN:6 23.505 
R237 ZN:6 ZN:4 0.56876 
R238 M6:DRN ZN:4 14.9999 
R239 M8:DRN ZN:4 22.2995 
R240 M4:DRN ZN:4 15.3563 
R241 M2:DRN ZN:4 15.5398 
R242 ZN:4 M10:DRN 42.451 
R243 M10:DRN M9:SRC 0.001 
R244 ZN:5 M20:DRN 15.5479 
R245 M20:DRN M19:SRC 0.001 
R246 M33:SRC M34:DRN 0.001 
R247 ZN:5 M18:DRN 14.9999 
R248 M18:DRN M17:SRC 0.001 
R249 M1:SRC M2:DRN 0.001 
R250 M2:DRN M4:DRN 1300.69 
R251 M4:DRN M3:SRC 0.001 
R252 M38:DRN M37:SRC 0.001 
R253 M8:DRN M7:SRC 0.001 
R254 M12:DRN M11:SRC 0.001 
R255 M6:DRN M5:SRC 0.001 
C256 M22:DRN 0 4.5e-18
C257 M24:SRC 0 7.31e-18
C258 M42:DRN 0 7.85e-18
C259 M32:DRN 0 6.28e-18
C260 ZN:1 0 4.99e-18
C261 M40:DRN 0 7.91e-18
C262 ZN:7 0 5.7961e-16
C263 M46:DRN 0 6.68e-18
C264 M26:DRN 0 1.08e-17
C265 M30:DRN 0 7.06e-18
C266 M28:DRN 0 7.27e-18
C267 M44:DRN 0 6.48e-18
C268 M48:DRN 0 9.96e-18
C269 M16:DRN 0 4.5e-18
C270 M36:DRN 0 1.59e-17
C271 M14:DRN 0 9.43e-18
C272 ZN:6 0 5.6726e-16
C273 M10:DRN 0 4.51e-18
C274 M20:DRN 0 4.5e-18
C275 M34:DRN 0 6.22e-18
C276 M18:DRN 0 4.5e-18
C277 M2:DRN 0 7.63e-18
C278 M4:DRN 0 4.84e-18
C279 M38:DRN 0 1.581e-17
C280 ZN 0 5.4e-19
C281 ZN:5 0 3.6e-19
C282 M8:DRN 0 4.5e-18
C283 M12:DRN 0 1.051e-17
C284 M6:DRN 0 4.54e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
