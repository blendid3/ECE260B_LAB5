.SUBCKT INVD3 I ZN
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.9e-07  AD=8e-14  AS=3.9e-14  PD=1.19e-06  PS=5.9e-07  SA=7.25e-07  SB=2.05e-07  NRD=0.566  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.65e-07  SB=4.65e-07  NRD=4.183  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=8e-14  PD=5.9e-07  PS=1.19e-06  SA=2.05e-07  SB=7.25e-07  NRD=4.141  NRS=0.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=1.07e-13  AS=5.2e-14  PD=1.45e-06  PS=7.2e-07  SA=7.25e-07  SB=2.05e-07  NRD=0.488  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.65e-07  SB=4.65e-07  NRD=2.057  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=1.07e-13  PD=7.2e-07  PS=1.45e-06  SA=2.05e-07  SB=7.25e-07  NRD=2.057  NRS=0.569  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M2:SRC M3:DRN 0.001 
R1 M3:DRN ZN 15.3129 
CC38208 M3:DRN M2:GATE 8.67e-18
CC38206 M3:DRN M3:GATE 4.203e-17
CC38202 M3:DRN I 2.401e-17
CC38189 M3:DRN I:1 4.132e-17
R2 M6:DRN ZN 15.4196 
R3 M4:DRN ZN 15.8634 
R4 ZN M1:DRN 15.7731 
CC38197 ZN M4:GATE 5.99e-18
CC38194 ZN M5:GATE 4.81e-18
CC38193 ZN M6:GATE 5.26e-18
CC38191 ZN I:1 3.91e-18
CC38210 ZN M1:GATE 8.81e-18
CC38207 ZN M2:GATE 5.4e-18
CC38205 ZN M3:GATE 7.7e-18
CC38204 ZN I 5.276e-17
R5 M1:DRN M4:DRN 1076.53 
CC38212 M1:DRN M1:GATE 4.174e-17
CC38200 M1:DRN M4:GATE 8.07e-18
CC38199 M4:DRN M4:GATE 4.582e-17
CC38188 M4:DRN I:1 1.79e-18
R6 M6:DRN M5:SRC 0.001 
CC38195 M6:DRN M5:GATE 4.573e-17
CC38192 M6:DRN M6:GATE 4.598e-17
CC38187 M6:DRN I:1 1.647e-17
C7 M3:DRN 0 5.19e-18
C8 ZN 0 3.4349e-16
C9 M1:DRN 0 2.638e-17
C10 M4:DRN 0 2.935e-17
C11 M6:DRN 0 1.212e-17
R12 M1:GATE M4:GATE 635.948 
R13 M4:GATE I:1 164.389 
R14 M2:GATE I:1 94.0755 
R15 M5:GATE I:1 111.3 
R16 M1:GATE I:1 138.947 
R17 I I:1 85.1298 
R18 M3:GATE I:1 194.508 
R19 I:1 M6:GATE 230.123 
R20 I M6:GATE 389.635 
R21 M6:GATE M3:GATE 890.253 
R22 M3:GATE I 329.333 
C23 M4:GATE 0 9.946e-17
C24 I:1 0 1.0923e-16
C25 M6:GATE 0 7.995e-17
C26 M3:GATE 0 3.221e-17
C27 I 0 1.04e-16
C28 M1:GATE 0 2.687e-17
C29 M5:GATE 0 1.0133e-16
C30 M2:GATE 0 5.564e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
