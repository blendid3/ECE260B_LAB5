.SUBCKT XNR2D0 A1 A2 ZN
MMM10 M9:SRC M10:GATE M10:SRC vdd pch L=6e-08 W=2.65e-07  AD=3e-14  AS=3.7e-14  PD=5.7e-07  PS=6.58e-07  SA=2.11e-07  SB=3.16e-07  NRD=0.48  NRS=0.572  SCA=7.419  SCB=0.008  SCC=0.0002752 
MMM11 M10:SRC M11:GATE vdd vdd pch L=6e-08 W=2.16e-07  AD=3e-14  AS=3.7e-14  PD=5.32e-07  PS=7.06e-07  SA=1.5e-07  SB=3.14e-07  NRD=0.69  NRS=0.972  SCA=17.254  SCB=0.019  SCC=0.002 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=2.04e-07  AD=3.6e-14  AS=2.4e-14  PD=7.6e-07  PS=4.45e-07  SA=5.07e-07  SB=1.85e-07  NRD=0.996  NRS=0.844  SCA=15.959  SCB=0.019  SCC=0.002 
MMM12 vdd M12:GATE M12:SRC vdd pch L=6e-08 W=2.67e-07  AD=4.6e-14  AS=4.3e-14  PD=8.74e-07  PS=8.5e-07  SA=1.65e-07  SB=1.72e-07  NRD=0.869  NRS=0.72  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=2.09e-07  AD=2.4e-14  AS=3.3e-14  PD=4.45e-07  PS=6.1e-07  SA=1.89e-07  SB=4.95e-07  NRD=0.844  NRS=0.87  SCA=15.959  SCB=0.019  SCC=0.002 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=1.97e-07  AD=3.9e-14  AS=2e-14  PD=6.42e-07  PS=4e-07  SA=6.41e-07  SB=1.9e-07  NRD=1.077  NRS=5.331  SCA=18.359  SCB=0.02  SCC=0.002 
MMM4 M2:SRC M4:GATE M3:DRN vss nch L=6e-08 W=2.05e-07  AD=3.3e-14  AS=4e-14  PD=6.1e-07  PS=6.58e-07  SA=2.15e-07  SB=1.87e-07  NRD=0.87  NRS=1.05  SCA=5.916  SCB=0.006  SCC=9.071e-05 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=2.04e-07  AD=3.3e-14  AS=2.1e-14  PD=7.3e-07  PS=4.36e-07  SA=1.65e-07  SB=4.26e-07  NRD=0.881  NRS=6.127  SCA=14.564  SCB=0.017  SCC=0.001 
MMM6 M3:SRC M6:GATE vss vss nch L=6.2e-08 W=1.93e-07  AD=2e-14  AS=2e-14  PD=4e-07  PS=4.14e-07  SA=3.49e-07  SB=4.6e-07  NRD=5.331  NRS=2.997  SCA=18.359  SCB=0.02  SCC=0.002 
MMM7 M7:DRN M7:GATE vdd vdd pch L=6e-08 W=2.66e-07  AD=4.4e-14  AS=3.9e-14  PD=8.6e-07  PS=6.35e-07  SA=3.7e-07  SB=1.7e-07  NRD=0.737  NRS=0.78  SCA=6.877  SCB=0.008  SCC=0.0002134 
MMM8 vdd M8:GATE M8:SRC vdd pch L=6e-08 W=2.65e-07  AD=3.9e-14  AS=3.8e-14  PD=6.35e-07  PS=5.5e-07  SA=6.7e-07  SB=2.41e-07  NRD=0.78  NRS=0.582  SCA=15.255  SCB=0.017  SCC=0.002 
MMM9 M8:SRC M9:GATE M9:SRC vdd pch L=6e-08 W=2.63e-07  AD=3.8e-14  AS=3e-14  PD=5.5e-07  PS=5.7e-07  SA=2.47e-07  SB=6.32e-07  NRD=0.582  NRS=0.48  SCA=15.255  SCB=0.017  SCC=0.002 
R0 M7:DRN ZN 30.5658 
R1 ZN M1:DRN 30.2705 
CC29315 ZN M3:DRN 6.102e-17
CC29309 ZN M1:GATE 1.253e-17
CC29295 ZN M7:GATE 8.77e-18
CC29287 ZN A2 9.43e-18
CC29308 M1:DRN M1:GATE 3.189e-17
CC29301 M7:DRN M9:SRC 1.47e-18
CC29292 M7:DRN M7:GATE 2.979e-17
C2 ZN 0 8.777e-17
C3 M1:DRN 0 1.584e-17
C4 M7:DRN 0 2.51e-17
R5 M7:GATE M1:GATE 312.999 
R6 M9:SRC M1:GATE 265.181 
R7 M1:GATE M3:DRN 271.97 
CC29307 M1:GATE M2:GATE 2.56e-18
CC29325 M1:GATE M12:SRC 5.232e-17
R8 M7:GATE M3:DRN 372.646 
R9 M3:DRN M9:SRC 75.5533 
CC29384 M3:DRN M4:GATE 2.4e-18
CC29338 M3:DRN M3:GATE 3.74e-17
CC29331 M3:DRN M9:GATE 2.415e-17
CC29373 M3:DRN M5:GATE 8.75e-18
CC29323 M3:DRN M12:SRC 6.41e-18
CC29316 M3:DRN A2 4.455e-17
CC29313 M3:DRN M2:SRC 8.33e-18
CC29312 M3:DRN M3:SRC 1.9e-18
CC29311 M3:DRN M6:GATE 5.492e-17
CC29381 M3:DRN M4:GATE 1.252e-17
R10 M9:SRC M7:GATE 363.348 
CC29304 M9:SRC M2:GATE 4.25e-18
CC29319 M9:SRC M12:SRC 1.398e-17
CC29298 M9:SRC M10:SRC 5.804e-17
CC29299 M9:SRC M8:SRC 5.339e-17
CC29300 M9:SRC M8:GATE 1.881e-17
CC29303 M9:SRC M2:SRC 1.818e-17
CC29328 M9:SRC M9:GATE 1.766e-17
CC29335 M9:SRC M3:GATE 1.559e-17
CC29350 M9:SRC M10:GATE 3.486e-17
CC29378 M9:SRC M4:GATE 2.18e-18
CC29360 M9:SRC A1 1.78e-18
CC29291 M7:GATE M8:GATE 4.71e-18
CC29296 M7:GATE A2 5.31e-18
C11 M1:GATE 0 2.289e-17
C12 M3:DRN 0 1.057e-17
C13 M9:SRC 0 2.605e-17
C14 M7:GATE 0 8.306e-17
R15 M2:GATE M8:GATE 300.147 
R16 M8:GATE A2 115.236 
CC29279 M8:GATE M8:SRC 1.184e-17
CC29280 M8:GATE M2:SRC 4.63e-18
R17 A2 M2:GATE 98.0127 
CC29282 A2 M8:SRC 8.65e-18
CC29283 A2 M2:SRC 7.432e-17
CC29285 M2:GATE M2:SRC 1.985e-17
C18 M8:GATE 0 4.211e-17
C19 A2 0 3.146e-17
C20 M2:GATE 0 3.358e-17
R21 M8:SRC M6:GATE 167.448 
R22 M2:SRC M6:GATE 163.888 
R23 M6:GATE M11:GATE 137.8 
CC29276 M6:GATE M3:SRC 2.647e-17
CC29362 M6:GATE A1 6.29e-18
CC29370 M6:GATE M5:GATE 9.99e-18
CC29273 M11:GATE M3:SRC 1.959e-17
CC29272 M11:GATE M10:SRC 3.519e-17
CC29367 M11:GATE M5:GATE 4.52e-18
CC29348 M11:GATE M10:GATE 1.77e-18
CC29342 M11:GATE M12:GATE 1.53e-18
CC29317 M11:GATE M12:SRC 4.39e-18
CC29326 M11:GATE M9:GATE 3.13e-18
CC29358 M11:GATE A1 1.212e-17
R24 M2:SRC M8:SRC 74.2419 
CC29382 M2:SRC M4:GATE 3.431e-17
CC29339 M2:SRC M3:GATE 1.473e-17
CC29277 M2:SRC M10:SRC 2.038e-17
CC29324 M2:SRC M12:SRC 3.09e-18
CC29278 M2:SRC M3:SRC 1.85e-18
CC29374 M2:SRC M5:GATE 5.73e-18
CC29329 M8:SRC M9:GATE 1.874e-17
CC29320 M8:SRC M12:SRC 2.63e-18
C25 M6:GATE 0 3.783e-17
C26 M11:GATE 0 4.049e-17
C27 M2:SRC 0 1.169e-17
C28 M8:SRC 0 1.2081e-16
R29 M10:SRC M3:SRC 60.4296 
CC29327 M10:SRC M9:GATE 6.77e-18
CC29318 M10:SRC M12:SRC 4.36e-18
CC29359 M10:SRC A1 1.23e-18
CC29349 M10:SRC M10:GATE 2.376e-17
CC29343 M10:SRC M12:GATE 3.27e-18
CC29337 M3:SRC M3:GATE 2.733e-17
CC29322 M3:SRC M12:SRC 2.842e-17
CC29363 M3:SRC A1 2.612e-17
CC29354 M3:SRC M10:GATE 3.91e-18
CC29371 M3:SRC M5:GATE 2.8e-18
C30 M10:SRC 0 8.34e-18
C31 M3:SRC 0 1.765e-17
R32 M4:GATE M5:GATE 385.045 
R33 M12:GATE M5:GATE 585.923 
R34 M5:GATE A1 99.9997 
CC29372 M5:GATE M5:DRN 2.899e-17
CC29366 M5:GATE M12:SRC 1.44e-17
CC29375 M5:GATE M3:GATE 2.92e-18
R35 A1 M12:GATE 193.466 
CC29364 A1 M5:DRN 6.978e-17
CC29357 A1 M12:SRC 7.55e-18
R36 M12:GATE M10:GATE 314.025 
CC29341 M12:GATE M12:SRC 2.661e-17
CC29351 M10:GATE M9:GATE 5.48e-18
CC29347 M10:GATE M12:SRC 1.219e-17
CC29383 M4:GATE M3:GATE 1.1e-18
C37 M5:GATE 0 1.3654e-16
C38 A1 0 7.259e-17
C39 M12:GATE 0 1.2967e-16
C40 M10:GATE 0 3.589e-17
C41 M4:GATE 0 6.03e-17
R42 M3:GATE M9:GATE 209.349 
R43 M12:SRC M9:GATE 213.369 
R44 M9:GATE M5:DRN 220.757 
R45 M5:DRN M12:SRC 71.0255 
C46 M3:GATE 0 1.47e-17
C47 M9:GATE 0 8.536e-17
C48 M5:DRN 0 1.2551e-16
C49 M12:SRC 0 5.41e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
