.SUBCKT OR2D0 A1 A2 Z
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=2.04e-07  AD=3.4e-14  AS=2.4e-14  PD=7.4e-07  PS=4.45e-07  SA=7.8e-07  SB=1.75e-07  NRD=0.947  NRS=0.844  SCA=18.109  SCB=0.02  SCC=0.002 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=2.04e-07  AD=2.4e-14  AS=2e-14  PD=4.45e-07  PS=4.05e-07  SA=4.7e-07  SB=4.85e-07  NRD=0.844  NRS=5.196  SCA=18.109  SCB=0.02  SCC=0.002 
MMM3 M2:SRC M3:GATE vss vss nch L=6e-08 W=2.04e-07  AD=2e-14  AS=3.9e-14  PD=4.05e-07  PS=7.9e-07  SA=2e-07  SB=7.55e-07  NRD=5.196  NRS=1.534  SCA=18.109  SCB=0.02  SCC=0.002 
MMM4 M4:DRN M4:GATE vdd vdd pch L=6e-08 W=2.63e-07  AD=4.5e-14  AS=3.6e-14  PD=8.7e-07  PS=5.4e-07  SA=7.75e-07  SB=1.75e-07  NRD=0.754  NRS=0.759  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=2.64e-07  AD=3.6e-14  AS=2.6e-14  PD=5.4e-07  PS=4.6e-07  SA=4.35e-07  SB=5.15e-07  NRD=0.759  NRS=4.018  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM6 M5:SRC M6:GATE M6:SRC vdd pch L=6e-08 W=2.6e-07  AD=2.6e-14  AS=4.5e-14  PD=4.6e-07  PS=8.7e-07  SA=1.75e-07  SB=7.75e-07  NRD=4.018  NRS=0.754  SCA=4.031  SCB=0.003  SCC=2.015e-05 
R0 M1:DRN Z 30.2324 
R1 Z M4:DRN 30.6659 
CC10184 Z M6:SRC 8.215e-17
CC10186 Z M1:GATE 3.78e-18
CC10183 Z M4:GATE 1.358e-17
CC10182 M4:DRN M4:GATE 2.945e-17
CC10188 M1:DRN M2:SRC 2.71e-17
CC10185 M1:DRN M1:GATE 5.7e-18
C2 Z 0 8.148e-17
C3 M4:DRN 0 2.529e-17
C4 M1:DRN 0 1.56e-17
R5 M4:GATE M1:GATE 371.924 
R6 M6:SRC M1:GATE 213.972 
R7 M1:GATE M2:SRC 211.407 
CC10196 M1:GATE A2 2.441e-17
CC10208 M1:GATE A1 3.183e-17
R8 M4:GATE M2:SRC 518.048 
R9 M2:SRC M6:SRC 78.0475 
CC10202 M2:SRC M6:GATE 4.54e-18
CC10192 M2:SRC M5:GATE 7.34e-18
CC10197 M2:SRC M2:GATE 2.169e-17
CC10195 M2:SRC A2 5.175e-17
CC10210 M2:SRC M3:GATE 2.044e-17
CC10206 M2:SRC A1 1.826e-17
R10 M6:SRC M4:GATE 524.334 
CC10204 M6:SRC A1 4.54e-18
CC10199 M6:SRC M6:GATE 2.986e-17
CC10193 M6:SRC A2 6.007e-17
CC10191 M4:GATE M5:GATE 8.61e-18
C11 M1:GATE 0 5.932e-17
C12 M2:SRC 0 9.417e-17
C13 M6:SRC 0 4.983e-17
C14 M4:GATE 0 8.151e-17
R15 M5:GATE M2:GATE 503.875 
R16 M2:GATE A2 84.5081 
CC10211 M2:GATE M3:GATE 1.86e-18
CC10207 M2:GATE A1 1.18e-17
R17 A2 M5:GATE 207.086 
CC10203 A2 M6:GATE 5.67e-18
CC10209 A2 A1 3.292e-17
CC10200 M5:GATE M6:GATE 1.998e-17
C18 M2:GATE 0 2.561e-17
C19 A2 0 1.114e-17
C20 M5:GATE 0 6.887e-17
R21 M3:GATE A1 83.4241 
R22 A1 M6:GATE 207.187 
R23 M6:GATE M3:GATE 489.272 
C24 A1 0 5.939e-17
C25 M6:GATE 0 4.583e-17
C26 M3:GATE 0 3.405e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
