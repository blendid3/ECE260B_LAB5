.SUBCKT MUX2D2 I0 I1 S Z
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=2.67e-07  AD=4.3e-14  AS=4.9e-14  PD=8.5e-07  PS=6.8e-07  SA=1.65e-07  SB=2.85e-07  NRD=0.72  NRS=0.867  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM11 M8:DRN M11:GATE M9:SRC vdd pch L=6e-08 W=4.15e-07  AD=4.6e-14  AS=5.8e-14  PD=7.98e-07  PS=8.42e-07  SA=2.81e-07  SB=2.7e-07  NRD=0.395  NRS=0.398  SCA=5.422  SCB=0.005  SCC=0.0001255 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7.4e-14  AS=3.9e-14  PD=1.16e-06  PS=5.9e-07  SA=9.08e-07  SB=1.9e-07  NRD=0.619  NRS=4.141  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM12 vdd M12:GATE M12:SRC vdd pch L=6e-08 W=5.24e-07  AD=6.8e-14  AS=5.2e-14  PD=1.3e-06  PS=7.2e-07  SA=9.64e-07  SB=1.3e-07  NRD=1.865  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=4.5e-14  PD=5.9e-07  PS=6.2e-07  SA=6.25e-07  SB=4.5e-07  NRD=4.141  NRS=0.349  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM13 M13:DRN M13:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=6.51e-07  SB=3.9e-07  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=4.5e-14  AS=4.8e-14  PD=6.2e-07  PS=7.61e-07  SA=2.85e-07  SB=7.4e-07  NRD=0.349  NRS=4.244  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM14 M8:SRC M14:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=6.6e-14  AS=4.7e-14  PD=9.2e-07  PS=7e-07  SA=3.1e-07  SB=6.3e-07  NRD=0.327  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE M4:SRC vss nch L=6e-08 W=2.33e-07  AD=3.3e-14  AS=2.3e-14  PD=6.26e-07  PS=4.3e-07  SA=6.33e-07  SB=2.33e-07  NRD=0.639  NRS=7.015  SCA=16.543  SCB=0.019  SCC=0.002 
MMM5 M3:SRC M5:GATE M4:DRN vss nch L=6e-08 W=2.51e-07  AD=3e-14  AS=3.4e-14  PD=4.69e-07  PS=6.54e-07  SA=1.73e-07  SB=1.025e-06  NRD=0.535  NRS=0.616  SCA=5.995  SCB=0.006  SCC=0.0001062 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=1.99e-07  AD=3.5e-14  AS=2e-14  PD=7.5e-07  PS=3.95e-07  SA=1.8e-07  SB=8.63e-07  NRD=0.972  NRS=0.553  SCA=13.679  SCB=0.016  SCC=0.001 
MMM7 M4:SRC M7:GATE vss vss nch L=6e-08 W=2.3e-07  AD=2.3e-14  AS=2.4e-14  PD=4.3e-07  PS=4.65e-07  SA=3.47e-07  SB=5.41e-07  NRD=7.015  NRS=9.028  SCA=16.543  SCB=0.019  SCC=0.002 
MMM8 M8:DRN M8:GATE M8:SRC vdd pch L=6e-08 W=3.53e-07  AD=3.9e-14  AS=4.4e-14  PD=6.82e-07  PS=6.2e-07  SA=2.96e-07  SB=9.4e-07  NRD=0.366  NRS=0.395  SCA=12.653  SCB=0.014  SCC=0.001 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=3.47e-07  AD=6.4e-14  AS=4.8e-14  PD=8.9e-07  PS=6.98e-07  SA=2.5e-07  SB=4.19e-07  NRD=0.78  NRS=0.452  SCA=12.895  SCB=0.014  SCC=0.001 
R0 M7:GATE I0 108.917 
R1 I0 M9:GATE 115.472 
CC3033 I0 M4:SRC 6.418e-17
CC3030 I0 M9:SRC 5.72e-18
CC3078 I0 M10:GATE 2.72e-18
CC3085 I0 S 5.49e-17
CC3094 I0 M6:GATE 4.2e-18
CC3043 I0 M8:GATE 6.06e-18
CC3038 I0 M10:DRN 1.587e-17
R2 M9:GATE M7:GATE 345.689 
CC3031 M9:GATE M4:SRC 1.7e-18
CC3036 M9:GATE M10:DRN 5.49e-18
CC3028 M9:GATE M9:SRC 3.518e-17
CC3071 M9:GATE M11:GATE 3.34e-18
CC3075 M9:GATE M10:GATE 2.78e-18
CC3081 M9:GATE S 1.358e-17
CC3032 M7:GATE M4:SRC 2.916e-17
CC3029 M7:GATE M9:SRC 3.89e-18
CC3089 M7:GATE M6:GATE 5.06e-18
CC3046 M7:GATE M4:GATE 1.76e-18
CC3040 M7:GATE M8:GATE 2.8e-18
C3 I0 0 3.651e-17
C4 M9:GATE 0 3.643e-17
C5 M7:GATE 0 3.383e-17
R6 Z M12:SRC 30.6479 
R7 M12:SRC M13:DRN 0.001 
CC3103 M12:SRC N_9:1 5.35e-18
CC3117 M12:SRC M13:GATE 2.883e-17
CC3125 M12:SRC M12:GATE 3.113e-17
R8 Z M2:DRN 15.2978 
R9 M2:DRN M1:SRC 0.001 
CC3112 M2:DRN N_9:1 8.901e-17
CC3062 M2:DRN I1 1.02e-18
CC3151 M2:DRN M2:GATE 1.378e-17
CC3146 M2:DRN M1:GATE 7.92e-18
CC3113 Z N_9:1 1.252e-17
CC3063 Z I1 1.359e-17
CC3163 Z M4:DRN 5.93e-17
CC3148 Z M2:GATE 3.27e-18
CC3144 Z M1:GATE 1.668e-17
CC3127 Z M12:GATE 3.151e-17
CC3122 Z M13:GATE 6.44e-18
C10 M12:SRC 0 7.56e-18
C11 M2:DRN 0 7.95e-18
C12 Z 0 1.0715e-16
R13 M4:GATE M8:GATE 247.775 
CC3045 M4:GATE M9:SRC 1.77e-18
CC3048 M4:GATE M4:SRC 2.761e-17
CC3093 M4:GATE M6:GATE 3.55e-18
CC3100 M4:GATE M5:GATE 1.34e-18
CC3139 M4:GATE M8:DRN 2.07e-18
CC3044 M4:GATE M8:SRC 3.405e-17
CC3110 M4:GATE N_9:1 1.78e-18
CC3162 M4:GATE M4:DRN 3.346e-17
CC3061 M4:GATE I1 7.63e-18
R14 M6:DRN M8:GATE 222.279 
R15 M8:GATE M10:DRN 214.198 
CC3106 M8:GATE N_9:1 4.65e-17
CC3096 M8:GATE M5:GATE 3.29e-18
CC3039 M8:GATE M9:SRC 1.28e-17
CC3135 M8:GATE M8:DRN 3.289e-17
CC3041 M8:GATE M3:SRC 4.12e-18
CC3140 M8:GATE M4:DRN 1.29e-18
CC3042 M8:GATE M4:SRC 2.21e-18
CC3157 M8:GATE M4:DRN 8.7e-18
CC3072 M8:GATE M11:GATE 5.12e-18
CC3054 M8:GATE M14:GATE 4.66e-18
R16 M10:DRN M6:DRN 71.088 
CC3087 M10:DRN M6:GATE 1.524e-17
CC3134 M10:DRN M8:DRN 2.609e-17
CC3035 M10:DRN M9:SRC 3.906e-17
CC3034 M10:DRN M8:SRC 1.096e-17
CC3156 M10:DRN M4:DRN 1.565e-17
CC3074 M10:DRN M10:GATE 3.218e-17
CC3070 M10:DRN M11:GATE 1.277e-17
CC3053 M10:DRN M14:GATE 1.44e-18
CC3080 M10:DRN S 2.09e-18
CC3084 M6:DRN S 7.802e-17
CC3090 M6:DRN M6:GATE 2.361e-17
C17 M4:GATE 0 1.288e-17
C18 M8:GATE 0 5.705e-17
C19 M10:DRN 0 7.081e-17
C20 M6:DRN 0 1.359e-16
R21 M11:GATE M10:GATE 307.4 
CC3132 M11:GATE M8:DRN 3.191e-17
CC3105 M11:GATE N_9:1 3.8e-18
CC3069 M11:GATE M9:SRC 2.54e-17
R22 M6:GATE M10:GATE 604.649 
R23 M10:GATE S 190.278 
CC3073 M10:GATE M9:SRC 6.52e-18
R24 S M6:GATE 104.357 
CC3079 S M9:SRC 2.68e-18
R25 M6:GATE M5:GATE 378.418 
CC3158 M6:GATE M4:DRN 8.3e-18
CC3107 M6:GATE N_9:1 1.41e-18
CC3086 M6:GATE M9:SRC 1.39e-18
CC3092 M6:GATE M4:SRC 5.09e-18
CC3143 M5:GATE M4:DRN 2.35e-18
CC3159 M5:GATE M4:DRN 1.937e-17
CC3108 M5:GATE N_9:1 3.37e-18
CC3095 M5:GATE M8:SRC 6.82e-18
CC3098 M5:GATE M3:SRC 3.446e-17
C26 M11:GATE 0 3.442e-17
C27 M10:GATE 0 1.2852e-16
C28 S 0 5.114e-17
C29 M6:GATE 0 1.3915e-16
C30 M5:GATE 0 6.024e-17
R31 M9:SRC M4:SRC 60.9906 
CC3104 M9:SRC N_9:1 2.784e-17
CC3131 M9:SRC M8:DRN 1.37e-18
CC3153 M9:SRC M4:DRN 2.1e-18
CC3138 M4:SRC M8:DRN 5.658e-17
C32 M9:SRC 0 2.431e-17
C33 M4:SRC 0 6.57e-18
R34 M8:SRC M3:SRC 60.9052 
CC3058 M8:SRC I1 5.897e-17
CC3051 M8:SRC M14:GATE 1.532e-17
CC3064 M8:SRC M3:GATE 6.62e-18
CC3152 M8:SRC M4:DRN 1.92e-18
CC3130 M8:SRC M8:DRN 1.88e-18
CC3102 M8:SRC N_9:1 5.032e-17
CC3055 M3:SRC M14:GATE 1.94e-18
CC3060 M3:SRC I1 2.168e-17
CC3065 M3:SRC M3:GATE 2.88e-18
CC3137 M3:SRC M8:DRN 6.582e-17
C35 M8:SRC 0 7.38e-18
C36 M3:SRC 0 3.982e-17
R37 M14:GATE M3:GATE 555.472 
R38 M3:GATE I1 129.901 
CC3111 M3:GATE N_9:1 2.46e-18
CC3149 M3:GATE M2:GATE 3.03e-18
R39 I1 M14:GATE 139.742 
CC3123 I1 M13:GATE 1.72e-18
CC3114 I1 N_9:1 2.02e-18
CC3164 I1 M4:DRN 4.257e-17
CC3147 I1 M2:GATE 2.32e-18
CC3128 I1 M12:GATE 2.27e-18
CC3101 M14:GATE N_9:1 2.334e-17
CC3115 M14:GATE M13:GATE 1.502e-17
C40 M3:GATE 0 5.556e-17
C41 I1 0 5.104e-17
C42 M14:GATE 0 5.197e-17
R43 N_9:1 M8:DRN 76.7473 
R44 M8:DRN M4:DRN 100.177 
R45 M4:DRN N_9:1 79.3539 
R46 M2:GATE N_9:1 91.2522 
R47 M13:GATE N_9:1 108.651 
R48 M12:GATE N_9:1 157.319 
R49 N_9:1 M1:GATE 147.727 
R50 M1:GATE M12:GATE 680.99 
C51 M8:DRN 0 2.87e-18
C52 M4:DRN 0 2.162e-17
C53 N_9:1 0 5.794e-17
C54 M1:GATE 0 6.046e-17
C55 M12:GATE 0 5.433e-17
C56 M13:GATE 0 3.889e-17
C57 M2:GATE 0 4.046e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
