.SUBCKT BUFFD4 I Z
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=6.7e-07  SB=9.3e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=4.3e-07  SB=1.17e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.6e-14  AS=3.9e-14  PD=1.12e-06  PS=5.9e-07  SA=1.43e-06  SB=1.7e-07  NRD=0.485  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M11:SRC M12:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.8e-14  PD=7.2e-07  PS=1.38e-06  SA=1.7e-07  SB=1.43e-06  NRD=2.057  NRS=0.538  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=1.17e-06  SB=4.3e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=9.3e-07  SB=6.7e-07  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=6.7e-07  SB=9.3e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=4.3e-07  SB=1.17e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M5:SRC M6:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.6e-14  PD=5.9e-07  PS=1.12e-06  SA=1.7e-07  SB=1.43e-06  NRD=4.141  NRS=0.583  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vdd M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.8e-14  AS=5.2e-14  PD=1.38e-06  PS=7.2e-07  SA=1.43e-06  SB=1.7e-07  NRD=0.44  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.17e-06  SB=4.3e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=9.3e-07  SB=6.7e-07  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M7:SRC M8:DRN 0.001 
R1 Z M8:DRN 15.3342 
R2 M8:DRN M10:DRN 1726.93 
CC77863 M8:DRN M8:GATE 4.59e-17
CC77864 M8:DRN M7:GATE 4.576e-17
CC77839 M8:DRN N_15:1 1.294e-17
CC77847 M8:DRN N_15:2 3.19e-18
R3 Z M10:DRN 15.6362 
R4 M10:DRN M9:SRC 0.001 
CC77887 M10:DRN M5:SRC 1.72e-18
CC77838 M10:DRN N_15:1 1.646e-17
CC77853 M10:DRN M10:GATE 4.619e-17
CC77857 M10:DRN M9:GATE 4.609e-17
R5 Z M2:DRN 15.3066 
R6 M2:DRN M1:SRC 0.001 
CC77874 M2:DRN M2:GATE 8.26e-18
CC77876 M2:DRN M1:GATE 2.132e-17
CC77842 M2:DRN N_15:1 1.495e-17
CC77849 M2:DRN N_15:2 6.924e-17
R7 Z M4:DRN 15.5544 
CC77866 Z M7:GATE 5.87e-18
CC77869 Z M11:SRC 1.9e-18
CC77872 Z M2:GATE 8.16e-18
CC77875 Z M1:GATE 2.82e-18
CC77880 Z M3:GATE 7.57e-18
CC77843 Z N_15:1 1.1495e-16
CC77850 Z N_15:2 7.19e-18
CC77854 Z M10:GATE 5e-18
CC77859 Z M9:GATE 1.199e-17
CC77861 Z M8:GATE 1.264e-17
CC77891 Z M5:SRC 1.706e-17
R8 M4:DRN M3:SRC 0.001 
CC77878 M4:DRN M3:GATE 8.59e-18
CC77884 M4:DRN M4:GATE 8.25e-18
CC77890 M4:DRN M5:SRC 1.94e-18
CC77841 M4:DRN N_15:1 8.699e-17
CC77848 M4:DRN N_15:2 1.183e-17
C9 M8:DRN 0 7.9e-18
C10 M10:DRN 0 8.82e-18
C11 M2:DRN 0 7.48e-18
C12 Z 0 2.076e-16
C13 M4:DRN 0 8.25e-18
R14 M6:GATE I:1 94.0755 
R15 M12:GATE I:1 111.3 
R16 M11:GATE I:1 239.272 
R17 M5:GATE I:1 202.244 
R18 I:1 I 38.8497 
CC77871 I:1 M11:SRC 1.632e-17
CC77893 I:1 M5:SRC 5.74e-17
CC77845 I:1 N_15:1 7.06e-18
CC77855 I:1 M10:GATE 1.33e-18
R19 M11:GATE I 440.438 
R20 I M5:GATE 372.274 
CC77870 I M11:SRC 8.179e-17
CC77892 I M5:SRC 2.184e-17
CC77844 I N_15:1 7.79e-18
R21 M5:GATE M11:GATE 727.924 
CC77889 M5:GATE M5:SRC 1.321e-17
CC77882 M5:GATE M4:GATE 8.67e-18
CC77868 M11:GATE M11:SRC 4.599e-17
CC77886 M11:GATE M5:SRC 9.62e-18
CC77852 M11:GATE M10:GATE 1.522e-17
CC77867 M12:GATE M11:SRC 4.6e-17
CC77885 M12:GATE M5:SRC 4.56e-18
CC77888 M6:GATE M5:SRC 4.26e-17
C22 I:1 0 4.611e-17
C23 I 0 5.52e-17
C24 M5:GATE 0 5.08e-17
C25 M11:GATE 0 6.054e-17
C26 M12:GATE 0 7.602e-17
C27 M6:GATE 0 2.299e-17
R28 M3:GATE M9:GATE 1165 
R29 N_15:2 M9:GATE 277.978 
R30 M9:GATE N_15:1 262.921 
R31 M4:GATE N_15:1 82.3623 
R32 M3:GATE N_15:1 222.23 
R33 M10:GATE N_15:1 111.3 
R34 N_15:2 N_15:1 53.0259 
R35 M11:SRC N_15:1 60.3125 
R36 N_15:1 M5:SRC 60.0651 
R37 M5:SRC M11:SRC 42.8918 
R38 M2:GATE N_15:2 94.0755 
R39 M3:GATE N_15:2 234.957 
R40 M8:GATE N_15:2 111.3 
R41 M1:GATE N_15:2 138.947 
R42 N_15:2 M7:GATE 164.389 
R43 M7:GATE M1:GATE 635.948 
C44 M9:GATE 0 4.661e-17
C45 N_15:1 0 1.727e-17
C46 M5:SRC 0 7.98e-17
C47 M11:SRC 0 5.545e-17
C48 N_15:2 0 2.512e-17
C49 M7:GATE 0 9.81e-17
C50 M1:GATE 0 6.118e-17
C51 M8:GATE 0 5.733e-17
C52 M10:GATE 0 3.958e-17
C53 M3:GATE 0 3.882e-17
C54 M2:GATE 0 4.147e-17
C55 M4:GATE 0 3.224e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
