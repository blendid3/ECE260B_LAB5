.SUBCKT OAI21D0 A1 A2 B ZN
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=2.01e-07  AD=2e-14  AS=2.4e-14  PD=3.95e-07  PS=4.45e-07  SA=4.85e-07  SB=4.6e-07  NRD=8.262  NRS=0.844  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM2 vss M2:GATE M1:DRN vss nch L=6e-08 W=2.02e-07  AD=3.9e-14  AS=2e-14  PD=7.9e-07  PS=3.95e-07  SA=7.45e-07  SB=2e-07  NRD=1.534  NRS=8.262  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM3 M3:DRN M3:GATE M1:SRC vss nch L=6e-08 W=2.01e-07  AD=3.4e-14  AS=2.4e-14  PD=7.4e-07  PS=4.45e-07  SA=1.75e-07  SB=7.7e-07  NRD=0.947  NRS=0.844  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM4 M4:DRN M4:GATE M4:SRC vdd pch L=6e-08 W=2.6e-07  AD=2.6e-14  AS=2.7e-14  PD=4.6e-07  PS=4.7e-07  SA=4.3e-07  SB=4.6e-07  NRD=4.054  NRS=0.404  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM5 M5:DRN M5:GATE vdd vdd pch L=6e-08 W=2.64e-07  AD=2.6e-14  AS=5.2e-14  PD=4.6e-07  PS=9.2e-07  SA=6.9e-07  SB=2e-07  NRD=4.054  NRS=1.386  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM6 M4:SRC M6:GATE vdd vdd pch L=6e-08 W=2.6e-07  AD=2.7e-14  AS=4.2e-14  PD=4.7e-07  PS=8.4e-07  SA=1.6e-07  SB=7.3e-07  NRD=0.404  NRS=0.704  SCA=4.031  SCB=0.003  SCC=2.015e-05 
R0 M3:DRN M1:DRN 60.7854 
CC92579 M3:DRN M1:SRC 3.63e-18
CC92577 M3:DRN ZN:1 3.14e-18
CC92598 M3:DRN A1 1.82e-18
CC92615 M3:DRN A2 3.298e-17
CC92604 M3:DRN M1:GATE 1.64e-18
CC92619 M3:DRN M3:GATE 2.856e-17
CC92576 M1:DRN ZN 7.411e-17
CC92585 M1:DRN B 1.042e-17
CC92589 M1:DRN M2:GATE 2.747e-17
CC92599 M1:DRN A1 5.04e-18
CC92605 M1:DRN M1:GATE 3.052e-17
C1 M3:DRN 0 8.519e-17
C2 M1:DRN 0 2.65e-17
R3 M4:GATE M1:GATE 854.594 
R4 M1:GATE A1 140.956 
CC92609 M1:GATE ZN:1 2.101e-17
CC92608 M1:GATE B 1.71e-18
CC92607 M1:GATE ZN 1.08e-18
CC92606 M1:GATE M2:GATE 1.38e-18
CC92621 M1:GATE M3:GATE 4.01e-18
R5 A1 M4:GATE 184.119 
CC92600 A1 M2:GATE 1.278e-17
CC92601 A1 ZN 4.047e-17
CC92602 A1 B 5.311e-17
CC92603 A1 ZN:1 1.452e-17
CC92595 A1 M5:GATE 2.84e-18
CC92596 A1 M5:DRN 1.41e-18
CC92622 A1 M3:GATE 1.22e-18
CC92613 A1 M6:GATE 6.45e-18
CC92617 A1 A2 3.741e-17
CC92590 M4:GATE M5:GATE 7.93e-18
CC92591 M4:GATE M5:DRN 3.043e-17
CC92592 M4:GATE ZN 4.78e-18
CC92593 M4:GATE B 3.68e-18
CC92594 M4:GATE ZN:1 2.32e-18
CC92611 M4:GATE M6:GATE 1.717e-17
CC92614 M4:GATE A2 1.17e-18
C6 M1:GATE 0 1.641e-17
C7 A1 0 2.023e-17
C8 M4:GATE 0 4.366e-17
R9 M1:SRC ZN:1 18.793 
R10 ZN:1 ZN 31.1686 
CC92623 ZN:1 M3:GATE 6.73e-18
CC92587 ZN:1 B 1.36e-18
CC92618 ZN:1 A2 2.241e-17
R11 ZN M5:DRN 31.0231 
CC92588 ZN M2:GATE 2.3e-18
CC92582 ZN M5:GATE 1.229e-17
CC92612 ZN M6:GATE 1.7e-18
CC92616 ZN A2 1.252e-17
CC92586 ZN B 9.264e-17
R12 M5:DRN M4:DRN 0.001 
CC92580 M5:DRN M5:GATE 2.975e-17
CC92583 M5:DRN B 2.38e-18
C13 M1:SRC 0 7e-19
C14 ZN:1 0 4.58e-18
C15 ZN 0 1.5194e-16
C16 M5:DRN 0 8.2e-18
R17 B M5:GATE 186.128 
R18 M5:GATE M2:GATE 882.056 
R19 M2:GATE B 143.183 
C20 M5:GATE 0 7.11e-17
C21 M2:GATE 0 3.696e-17
C22 B 0 2.705e-17
R23 A2 M3:GATE 139.26 
R24 M3:GATE M6:GATE 833.977 
R25 M6:GATE A2 182.597 
C26 M3:GATE 0 2.999e-17
C27 M6:GATE 0 8.012e-17
C28 A2 0 4.754e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
