.SUBCKT ND2D3 A1 A2 ZN
MMM10 M10:DRN M10:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=9.2e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vdd M11:GATE M11:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=1.18e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.567  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=1.44e-06  NRD=2.099  NRS=0.532  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M1:SRC M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=1.18e-06  SB=4.2e-07  NRD=4.12  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=9.4e-07  SB=6.6e-07  NRD=7.648  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M3:SRC M4:GATE M4:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=9.2e-07  NRD=4.12  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 M5:DRN M5:GATE M5:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=1.18e-06  NRD=4.183  NRS=4.12  SCA=11.955  SCB=0.013  SCC=0.001 
MMM6 M5:SRC M6:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.2e-14  PD=5.9e-07  PS=1.1e-06  SA=1.6e-07  SB=1.44e-06  NRD=4.12  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vdd M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.44e-06  SB=1.6e-07  NRD=0.532  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.18e-06  SB=4.2e-07  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=9.4e-07  SB=6.6e-07  NRD=6.61  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
CC45059 M1:SRC A1 1.08e-18
CC45014 M5:SRC A2 1.08e-18
R0 M7:SRC ZN 29.9999 
R1 M4:SRC ZN 34.4232 
R2 M1:DRN ZN 33.1487 
R3 M9:SRC ZN 31.1674 
R4 ZN M11:SRC 31.9759 
CC45070 ZN M5:GATE 1.88e-18
CC45076 ZN M1:GATE 9.15e-18
CC45022 ZN M3:GATE 7.46e-18
CC45029 ZN A1:1 2.91e-18
CC45019 ZN M6:GATE 1.12e-18
CC45061 ZN A1 1.5993e-16
CC45003 ZN A2:1 1.354e-17
CC45049 ZN M7:GATE 1.862e-17
CC45011 ZN M8:GATE 1.193e-17
CC45036 ZN M11:GATE 4.46e-18
CC45008 ZN M9:GATE 7.08e-18
CC45016 ZN A2 1.1813e-16
CC45043 ZN M10:GATE 5.22e-18
CC45005 ZN M12:GATE 3.57e-18
CC45068 ZN M4:GATE 4.84e-18
CC45020 ZN M2:GATE 9.72e-18
R5 M9:SRC M11:SRC 1622.69 
R6 M11:SRC M12:DRN 0.001 
CC45004 M11:SRC M12:GATE 2.811e-17
CC45017 M11:SRC M6:GATE 1.9e-18
CC45012 M11:SRC A2 8.17e-18
CC45033 M11:SRC M11:GATE 2.809e-17
R7 M9:SRC M10:DRN 0.001 
CC45025 M9:SRC A1:1 1.39e-18
CC45013 M9:SRC A2 6.91e-18
CC45040 M9:SRC M10:GATE 2.867e-17
CC45006 M9:SRC M9:GATE 2.821e-17
R8 M1:DRN M4:SRC 643.825 
CC45060 M1:DRN A1 2.893e-17
R9 M4:SRC M5:DRN 0.001 
CC45073 M4:SRC M5:GATE 4.96e-18
CC45028 M4:SRC A1:1 3.309e-17
CC45056 M4:SRC A1 5.3e-18
CC45065 M4:SRC M4:GATE 2.891e-17
R10 M7:SRC M8:DRN 0.001 
CC45054 M7:SRC A1 5.53e-18
CC45048 M7:SRC M7:GATE 2.818e-17
CC45010 M7:SRC M8:GATE 2.775e-17
C11 ZN 0 2.1815e-16
C12 M11:SRC 0 1.281e-17
C13 M9:SRC 0 5.87e-18
C14 M1:DRN 0 3.143e-17
C15 M4:SRC 0 2.164e-17
C16 M7:SRC 0 3.89e-18
R17 M8:GATE A2 477.803 
R18 M2:GATE A2 403.857 
R19 A2:1 A2 39.4886 
R20 M12:GATE A2 144.989 
R21 A2 M6:GATE 123.225 
CC45030 A2 A1:1 1.169e-17
CC45075 A2 M1:GATE 6.89e-18
CC45037 A2 M11:GATE 6.58e-18
CC45044 A2 M10:GATE 6.35e-18
CC45062 A2 A1 1.2782e-16
CC45069 A2 M5:GATE 7.92e-18
R22 M6:GATE M12:GATE 543.896 
CC45027 M6:GATE A1:1 3.01e-18
CC45071 M6:GATE M5:GATE 4.14e-18
CC45023 M12:GATE A1:1 1.035e-17
CC45032 M12:GATE M11:GATE 7.66e-18
R23 M9:GATE A2:1 111.3 
CC45026 M9:GATE A1:1 1.85e-18
CC45041 M9:GATE M10:GATE 7.71e-18
R24 M3:GATE A2:1 94.0755 
R25 M8:GATE A2:1 223.959 
R26 A2:1 M2:GATE 189.298 
CC45074 A2:1 M1:GATE 1.095e-17
CC45031 A2:1 A1:1 6.46e-18
CC45045 A2:1 M10:GATE 3.19e-18
CC45063 A2:1 A1 9.25e-18
R27 M2:GATE M8:GATE 760.394 
CC45077 M2:GATE M1:GATE 3.82e-18
CC45058 M2:GATE A1 1.28e-17
CC45047 M8:GATE M7:GATE 7.78e-18
CC45057 M3:GATE A1 1.329e-17
CC45066 M3:GATE M4:GATE 3.95e-18
C28 A2 0 6.684e-17
C29 M6:GATE 0 5.545e-17
C30 M12:GATE 0 8.087e-17
C31 M9:GATE 0 5.042e-17
C32 A2:1 0 6.087e-17
C33 M2:GATE 0 2.855e-17
C34 M8:GATE 0 6.074e-17
C35 M3:GATE 0 2.264e-17
R36 A1 M1:GATE 124.765 
R37 M1:GATE M7:GATE 514.481 
R38 M7:GATE A1 151.23 
R39 M10:GATE A1 448.204 
R40 M4:GATE A1 378.839 
R41 A1 A1:1 37.7348 
R42 M5:GATE A1:1 94.0755 
R43 M10:GATE A1:1 238.184 
R44 M4:GATE A1:1 201.322 
R45 A1:1 M11:GATE 111.3 
R46 M4:GATE M10:GATE 722.167 
C47 M1:GATE 0 3.096e-17
C48 M7:GATE 0 8.493e-17
C49 A1 0 2.699e-17
C50 A1:1 0 2.965e-17
C51 M11:GATE 0 7.484e-17
C52 M4:GATE 0 2.292e-17
C53 M10:GATE 0 8.449e-17
C54 M5:GATE 0 3.162e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
