.SUBCKT AN2D1 A1 A2 Z
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=1.95e-07  AD=3.9e-14  AS=1.6e-14  PD=7.9e-07  PS=3.55e-07  SA=2e-07  SB=7.6e-07  NRD=1.069  NRS=20.501  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM2 M1:SRC M2:GATE vss vss nch L=6e-08 W=2.01e-07  AD=1.6e-14  AS=3.2e-14  PD=3.55e-07  PS=4.6e-07  SA=4.2e-07  SB=5.4e-07  NRD=20.501  NRS=0.956  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM3 M3:DRN M3:GATE vss vss nch L=6e-08 W=3.97e-07  AD=7e-14  AS=6.5e-14  PD=1.14e-06  PS=9.2e-07  SA=3.28e-07  SB=1.8e-07  NRD=0.6  NRS=0.761  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 vdd M4:GATE M4:SRC vdd pch L=6e-08 W=2.65e-07  AD=5.2e-14  AS=2.7e-14  PD=9.2e-07  PS=4.7e-07  SA=2e-07  SB=7.6e-07  NRD=0.84  NRS=0.438  SCA=6.553  SCB=0.007  SCC=0.00018 
MMM5 M4:SRC M5:GATE vdd vdd pch L=6e-08 W=2.68e-07  AD=2.7e-14  AS=3.9e-14  PD=4.7e-07  PS=5.13e-07  SA=4.7e-07  SB=4.9e-07  NRD=0.438  NRS=0.714  SCA=6.553  SCB=0.007  SCC=0.00018 
MMM6 M6:DRN M6:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=9.4e-14  AS=7.8e-14  PD=1.4e-06  PS=1.027e-06  SA=3.28e-07  SB=1.8e-07  NRD=0.453  NRS=0.755  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M6:DRN Z 15.4371 
R1 Z M3:DRN 30.4633 
CC75198 Z M1:DRN 8.815e-17
CC75193 Z M3:GATE 1.325e-17
CC75180 Z M6:GATE 5.04e-18
CC75191 M3:DRN M3:GATE 6.68e-18
CC75185 M3:DRN M4:SRC 2.209e-17
CC75182 M6:DRN M4:SRC 2.63e-18
CC75177 M6:DRN M6:GATE 4.511e-17
C2 Z 0 1.0343e-16
C3 M3:DRN 0 2.616e-17
C4 M6:DRN 0 3.247e-17
R5 M1:GATE A1 155.757 
R6 A1 M4:GATE 137.944 
CC75174 A1 M5:GATE 6.98e-18
CC75175 A1 A2 6.855e-17
CC75189 A1 M4:SRC 2.46e-18
CC75195 A1 M3:GATE 3.488e-17
CC75200 A1 M1:DRN 9.57e-18
R7 M4:GATE M1:GATE 682.92 
CC75173 M4:GATE A2 2.3e-18
CC75172 M4:GATE M5:GATE 8.02e-18
CC75184 M4:GATE M4:SRC 3.65e-17
CC75187 M1:GATE M4:SRC 4.78e-18
CC75197 M1:GATE M1:DRN 2.136e-17
CC75176 M1:GATE M2:GATE 4.82e-18
C8 A1 0 4.531e-17
C9 M4:GATE 0 5.158e-17
C10 M1:GATE 0 3.487e-17
R11 M2:GATE M5:GATE 682.92 
R12 M5:GATE A2 137.944 
CC75178 M5:GATE M6:GATE 3.41e-18
CC75183 M5:GATE M4:SRC 3.973e-17
R13 A2 M2:GATE 155.757 
CC75181 A2 M6:GATE 1.24e-17
CC75188 A2 M4:SRC 6.55e-18
CC75194 A2 M3:GATE 1.136e-17
CC75199 A2 M1:DRN 6.972e-17
CC75186 M2:GATE M4:SRC 1.536e-17
C14 M5:GATE 0 4.096e-17
C15 A2 0 2.625e-17
C16 M2:GATE 0 4.177e-17
R17 M1:DRN M3:GATE 309.393 
R18 M4:SRC M3:GATE 305.299 
R19 M3:GATE M6:GATE 388.973 
R20 M1:DRN M6:GATE 353.732 
R21 M6:GATE M4:SRC 349.055 
R22 M4:SRC M1:DRN 76.9717 
C23 M3:GATE 0 4.291e-17
C24 M6:GATE 0 1.0282e-16
C25 M4:SRC 0 1.29e-16
C26 M1:DRN 0 4.66e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
