.SUBCKT AN2D2 A1 A2 Z
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7.2e-14  AS=2.7e-14  PD=1.15e-06  PS=5.3e-07  SA=1.85e-07  SB=9.95e-07  NRD=0.609  NRS=13.316  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M1:SRC M2:GATE vss vss nch L=6.1e-08 W=3.93e-07  AD=2.7e-14  AS=5.8e-14  PD=5.3e-07  PS=6.9e-07  SA=3.85e-07  SB=7.95e-07  NRD=13.316  NRS=0.662  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.9e-07  AD=6.8e-14  AS=3.9e-14  PD=1.13e-06  PS=5.9e-07  SA=1.005e-06  SB=1.75e-07  NRD=0.592  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 vss M4:GATE M4:SRC vss nch L=6e-08 W=3.97e-07  AD=5.8e-14  AS=3.9e-14  PD=6.9e-07  PS=5.9e-07  SA=7.45e-07  SB=4.35e-07  NRD=0.662  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=5.24e-07  AD=1.04e-13  AS=5.5e-14  PD=1.44e-06  PS=7.3e-07  SA=2e-07  SB=9.8e-07  NRD=0.564  NRS=0.287  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M5:SRC M6:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.5e-14  AS=5.2e-14  PD=7.3e-07  PS=7.2e-07  SA=4.7e-07  SB=7.1e-07  NRD=0.287  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vdd M7:GATE M7:SRC vdd pch L=6e-08 W=5.2e-07  AD=9.6e-14  AS=5.3e-14  PD=1.41e-06  PS=7.25e-07  SA=9.95e-07  SB=1.85e-07  NRD=0.549  NRS=1.051  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 vdd M8:GATE M8:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.3e-14  PD=7.2e-07  PS=7.25e-07  SA=7.3e-07  SB=4.5e-07  NRD=2.099  NRS=1.051  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M1:GATE A1 124.451 
R1 A1 M5:GATE 142.288 
CC75570 A1 N_12:1 3.998e-17
CC75575 A1 M5:SRC 1.94e-18
CC75591 A1 M1:DRN 3.564e-17
CC75556 A1 M2:GATE 1.653e-17
CC75557 A1 A2 4.292e-17
R2 M5:GATE M1:GATE 538.172 
CC75564 M5:GATE N_12:1 2.01e-18
CC75572 M5:GATE M5:SRC 2.619e-17
CC75554 M5:GATE A2 2.02e-18
CC75553 M5:GATE M6:GATE 6.47e-18
CC75567 M1:GATE N_12:1 7.44e-18
CC75558 M1:GATE M2:GATE 5.65e-18
CC75559 M1:GATE A2 1.652e-17
C3 A1 0 3.629e-17
C4 M5:GATE 0 9.634e-17
C5 M1:GATE 0 2.765e-17
R6 M2:GATE M6:GATE 530.987 
R7 M6:GATE A2 155.219 
CC75563 M6:GATE N_12:1 2.071e-17
CC75571 M6:GATE M5:SRC 2.783e-17
CC75577 M6:GATE M8:GATE 6.47e-18
R8 A2 M2:GATE 113.322 
CC75569 A2 N_12:1 2.11e-18
CC75574 A2 M5:SRC 7.83e-17
CC75580 A2 M8:GATE 1.77e-18
CC75566 M2:GATE N_12:1 1.166e-17
C9 M6:GATE 0 8.467e-17
C10 A2 0 4.008e-17
C11 M2:GATE 0 2.476e-17
R12 M3:SRC M4:SRC 0.001 
R13 M4:SRC Z 15.2809 
CC75565 M4:SRC N_12:1 8.16e-17
CC75588 M4:SRC M3:GATE 2.607e-17
CC75586 M4:SRC M4:GATE 8.11e-18
R14 Z M8:SRC 15.4202 
CC75584 Z M4:GATE 2.94e-18
CC75573 Z M5:SRC 1.278e-17
CC75583 Z M7:GATE 2.051e-17
CC75579 Z M8:GATE 4.47e-18
CC75568 Z N_12:1 5.104e-17
CC75589 Z M1:DRN 3.869e-17
CC75587 Z M3:GATE 2.53e-18
R15 M8:SRC M7:SRC 0.001 
CC75562 M8:SRC N_12:1 6.69e-17
CC75581 M8:SRC M7:GATE 2.17e-18
CC75576 M8:SRC M8:GATE 4.31e-17
C16 M4:SRC 0 5.7e-18
C17 Z 0 1.4746e-16
C18 M8:SRC 0 9.42e-18
R19 M8:GATE N_12:1 104.675 
R20 M4:GATE N_12:1 93.1916 
R21 M3:GATE N_12:1 148.412 
R22 M7:GATE N_12:1 154.27 
R23 M5:SRC N_12:1 74.9033 
R24 N_12:1 M1:DRN 75.19 
R25 M1:DRN M5:SRC 105.906 
R26 M7:GATE M3:GATE 638.836 
C27 M8:GATE 0 7.271e-17
C28 N_12:1 0 7.958e-17
C29 M1:DRN 0 9.836e-17
C30 M5:SRC 0 3.415e-17
C31 M7:GATE 0 5.862e-17
C32 M3:GATE 0 6.443e-17
C33 M4:GATE 0 4.469e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
