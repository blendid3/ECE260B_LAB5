.SUBCKT NR2D1 A1 A2 ZN
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.6e-14  AS=3.9e-14  PD=1.12e-06  PS=5.9e-07  SA=4.3e-07  SB=1.7e-07  NRD=0.583  NRS=4.183  SCA=11.516  SCB=0.012  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=6.6e-14  AS=3.9e-14  PD=1.12e-06  PS=5.9e-07  SA=1.7e-07  SB=4.3e-07  NRD=0.583  NRS=4.183  SCA=11.516  SCB=0.012  SCC=0.001 
MMM3 M3:DRN M3:GATE M3:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.8e-14  AS=5.2e-14  PD=1.38e-06  PS=7.2e-07  SA=4.3e-07  SB=1.7e-07  NRD=0.538  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 vdd M4:GATE M3:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.8e-14  AS=5.2e-14  PD=1.38e-06  PS=7.2e-07  SA=1.7e-07  SB=4.3e-07  NRD=0.538  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M3:DRN ZN 30.5557 
R1 ZN M1:SRC 30.8974 
CC47614 ZN A1 7.736e-17
CC47613 ZN A2 9.2e-18
CC47612 ZN M1:GATE 1.535e-17
CC47611 ZN M2:GATE 5.01e-18
CC47610 ZN M3:GATE 7.27e-18
R2 M1:SRC M2:SRC 0.001 
CC47619 M1:SRC A1 2.596e-17
CC47618 M1:SRC A2 1.914e-17
CC47617 M1:SRC M1:GATE 6.49e-18
CC47616 M1:SRC M2:GATE 1.069e-17
CC47615 M1:SRC M3:GATE 1.43e-18
CC47608 M3:DRN A1 1.19e-18
CC47607 M3:DRN M3:GATE 2.845e-17
C3 ZN 0 1.5383e-16
C4 M1:SRC 0 9.25e-18
C5 M3:DRN 0 2.197e-17
R6 A1 M1:GATE 122.976 
R7 M1:GATE M3:GATE 550.193 
CC47603 M1:GATE M2:GATE 2.01e-18
R8 M3:GATE A1 146.667 
CC47599 M3:GATE M4:GATE 1.503e-17
CC47601 M3:GATE A2 1.389e-17
CC47600 A1 M4:GATE 2.48e-18
CC47602 A1 A2 2.423e-17
CC47604 A1 M2:GATE 8.57e-18
CC47605 A1 M3:SRC 1.05e-18
C9 M1:GATE 0 5.28e-17
C10 M3:GATE 0 4.082e-17
C11 A1 0 3.891e-17
R12 M2:GATE A2 119.055 
R13 A2 M4:GATE 143.093 
R14 M4:GATE M2:GATE 512.212 
C15 A2 0 1.0364e-16
C16 M4:GATE 0 1.0086e-16
C17 M2:GATE 0 4.637e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
