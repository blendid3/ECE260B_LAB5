.SUBCKT XNR2D1 A1 A2 ZN
MMM10 vdd M10:GATE M10:SRC vdd pch L=6e-08 W=2.64e-07  AD=4.5e-14  AS=4.2e-14  PD=7.45e-07  PS=8.4e-07  SA=1.6e-07  SB=1.75e-07  NRD=0.684  NRS=0.704  SCA=4.031  SCB=0.003  SCC=2.015e-05 
MMM11 M11:DRN M11:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=9.1e-14  AS=6.5e-14  PD=1.39e-06  PS=7.7e-07  SA=7.09e-07  SB=1.75e-07  NRD=0.541  NRS=0.66  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.8e-14  AS=4.9e-14  PD=1.13e-06  PS=6.4e-07  SA=5.87e-07  SB=1.75e-07  NRD=0.496  NRS=0.371  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M7:SRC M12:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.7e-14  AS=6.5e-14  PD=8.53e-07  PS=7.7e-07  SA=3.1e-07  SB=4.85e-07  NRD=4.762  NRS=0.66  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.97e-07  AD=4.9e-14  AS=4.2e-14  PD=6.4e-07  PS=7.48e-07  SA=2.3e-07  SB=4.85e-07  NRD=0.371  NRS=8.791  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE M3:SRC vss nch L=6e-08 W=1.95e-07  AD=3e-14  AS=1.9e-14  PD=5.63e-07  PS=3.9e-07  SA=6.26e-07  SB=1.99e-07  NRD=0.843  NRS=8.478  SCA=18.359  SCB=0.02  SCC=0.002 
MMM4 M2:SRC M4:GATE M3:DRN vss nch L=6e-08 W=2.36e-07  AD=2.4e-14  AS=3.6e-14  PD=4.32e-07  PS=6.67e-07  SA=1.74e-07  SB=7.45e-07  NRD=0.499  NRS=0.721  SCA=6.258  SCB=0.006  SCC=0.0001231 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=1.99e-07  AD=3.4e-14  AS=2.2e-14  PD=7.4e-07  PS=4.46e-07  SA=1.75e-07  SB=4.11e-07  NRD=0.947  NRS=1.704  SCA=13.679  SCB=0.016  SCC=0.001 
MMM6 M3:SRC M6:GATE vss vss nch L=6.2e-08 W=1.92e-07  AD=1.9e-14  AS=2.1e-14  PD=3.9e-07  PS=4.34e-07  SA=3.39e-07  SB=4.78e-07  NRD=8.478  NRS=0.609  SCA=18.359  SCB=0.02  SCC=0.002 
MMM7 M7:DRN M7:GATE M7:SRC vdd pch L=6e-08 W=3.72e-07  AD=3.9e-14  AS=4e-14  PD=6.97e-07  PS=6.07e-07  SA=2.64e-07  SB=7.55e-07  NRD=10.154  NRS=0.34  SCA=12.196  SCB=0.013  SCC=0.001 
MMM8 M7:DRN M8:GATE M8:SRC vdd pch L=6e-08 W=2.4e-07  AD=2.5e-14  AS=3.3e-14  PD=4.43e-07  PS=5.65e-07  SA=2.46e-07  SB=1.015e-06  NRD=0.476  NRS=0.612  SCA=6.833  SCB=0.007  SCC=0.000198 
MMM9 M8:SRC M9:GATE vdd vdd pch L=6e-08 W=2.66e-07  AD=3.6e-14  AS=4.5e-14  PD=6.25e-07  PS=7.45e-07  SA=1.7e-07  SB=3.16e-07  NRD=0.561  NRS=0.684  SCA=15.255  SCB=0.017  SCC=0.002 
R0 M3:SRC M8:SRC 60.6379 
CC29434 M3:SRC M3:DRN 7.156e-17
CC29401 M3:SRC M6:GATE 1.003e-17
CC29390 M3:SRC M3:GATE 3.081e-17
CC29398 M3:SRC M9:GATE 2.044e-17
CC29406 M3:SRC M2:SRC 3.043e-17
CC29494 M3:SRC M5:GATE 2.84e-18
CC29419 M8:SRC M7:DRN 2.26e-18
CC29389 M8:SRC M3:GATE 2.01e-18
CC29468 M8:SRC M10:GATE 3.46e-18
CC29385 M8:SRC M10:SRC 4.178e-17
CC29399 M8:SRC M6:GATE 4.87e-18
CC29396 M8:SRC M9:GATE 3.996e-17
CC29476 M8:SRC M8:GATE 2.36e-17
CC29387 M8:SRC M7:GATE 8.33e-18
CC29482 M8:SRC A1 2.255e-17
CC29431 M8:SRC M3:DRN 1.9e-18
C1 M3:SRC 0 6.44e-18
C2 M8:SRC 0 1.608e-17
R3 A1 M10:GATE 199.983 
R4 M8:GATE M10:GATE 317.206 
R5 M10:GATE M5:GATE 583.368 
CC29469 M10:GATE M7:DRN 2.28e-18
CC29467 M10:GATE M9:GATE 1.04e-18
CC29466 M10:GATE M10:SRC 2.93e-17
R6 A1 M5:GATE 96.8281 
R7 M5:GATE M4:GATE 383.19 
CC29497 M5:GATE M2:SRC 1.966e-17
CC29498 M5:GATE M3:GATE 2.87e-18
CC29489 M5:GATE M10:SRC 1.602e-17
CC29495 M5:GATE M5:DRN 3.108e-17
CC29500 M4:GATE M7:DRN 2.13e-18
CC29501 M4:GATE M7:GATE 3.35e-18
CC29504 M4:GATE M3:DRN 2.641e-17
CC29505 M4:GATE M2:SRC 4.606e-17
CC29506 M4:GATE M3:GATE 1.63e-18
CC29478 M8:GATE M7:GATE 5.95e-18
CC29477 M8:GATE M7:DRN 3.671e-17
CC29475 M8:GATE M9:GATE 3.26e-18
CC29474 M8:GATE M10:SRC 1.466e-17
CC29487 A1 M5:DRN 6.785e-17
CC29485 A1 M6:GATE 1.509e-17
CC29481 A1 M9:GATE 5.24e-18
CC29480 A1 M10:SRC 7.67e-18
C8 M10:GATE 0 1.2699e-16
C9 M5:GATE 0 1.3831e-16
C10 M4:GATE 0 5.183e-17
C11 M8:GATE 0 3.281e-17
C12 A1 0 7.397e-17
R13 M5:DRN M10:SRC 71.0738 
R14 M10:SRC M7:GATE 211.21 
CC29442 M10:SRC M12:GATE 2.63e-18
CC29430 M10:SRC M3:DRN 2.883e-17
CC29425 M10:SRC M1:GATE 6.55e-18
CC29417 M10:SRC M7:DRN 1.539e-17
CC29410 M10:SRC M11:GATE 1.148e-17
CC29404 M10:SRC M2:SRC 1.79e-18
CC29391 M10:SRC M7:SRC 5.61e-18
CC29395 M10:SRC M9:GATE 5.23e-18
R15 M3:GATE M7:GATE 230.551 
R16 M7:GATE M5:DRN 218.1 
CC29444 M7:GATE M12:GATE 3.24e-18
CC29432 M7:GATE M3:DRN 2.29e-17
CC29420 M7:GATE M7:DRN 2.185e-17
CC29405 M7:GATE M2:SRC 2.28e-18
CC29393 M7:GATE M7:SRC 2.343e-17
CC29400 M7:GATE M6:GATE 4.28e-18
CC29447 M3:GATE M12:GATE 2.33e-18
CC29436 M3:GATE M3:DRN 2.506e-17
CC29423 M3:GATE M7:DRN 2.868e-17
CC29407 M3:GATE M2:SRC 1.336e-17
CC29457 M3:GATE A2 4.96e-18
CC29394 M3:GATE M7:SRC 9.62e-18
C17 M10:SRC 0 5.477e-17
C18 M7:GATE 0 8.814e-17
C19 M5:DRN 0 1.3578e-16
C20 M3:GATE 0 1.138e-17
R21 M11:DRN ZN 30.6142 
R22 ZN M1:DRN 15.4687 
CC29460 ZN A2 1.44e-17
CC29414 ZN M11:GATE 1.662e-17
CC29428 ZN M1:GATE 1.102e-17
CC29438 ZN M3:DRN 5.717e-17
CC29413 M1:DRN M11:GATE 1.85e-18
CC29459 M1:DRN A2 1.11e-18
CC29427 M1:DRN M1:GATE 1.828e-17
CC29437 M1:DRN M3:DRN 3.506e-17
CC29409 M11:DRN M11:GATE 2.91e-17
CC29416 M11:DRN M7:DRN 3.11e-18
C23 ZN 0 1.142e-16
C24 M1:DRN 0 2.625e-17
C25 M11:DRN 0 3.161e-17
R26 M1:GATE M7:DRN 322.241 
R27 M11:GATE M7:DRN 336.935 
R28 M7:DRN M3:DRN 74.459 
CC29443 M7:DRN M12:GATE 1.375e-17
CC29462 M7:DRN M2:GATE 2.3e-18
CC29422 M7:DRN M2:SRC 6.73e-18
CC29421 M7:DRN M6:GATE 4.215e-17
CC29415 M7:DRN M7:SRC 7.607e-17
R29 M1:GATE M3:DRN 331.879 
R30 M3:DRN M11:GATE 347.009 
CC29435 M3:DRN M2:SRC 6.32e-18
CC29433 M3:DRN M6:GATE 1.4e-18
CC29455 M3:DRN A2 2.13e-18
R31 M11:GATE M1:GATE 382.107 
CC29440 M11:GATE M12:GATE 4.66e-18
CC29452 M11:GATE A2 6.52e-18
CC29458 M1:GATE A2 4.28e-17
CC29448 M1:GATE M12:GATE 2.96e-18
C32 M7:DRN 0 3.29e-17
C33 M3:DRN 0 5.25e-18
C34 M11:GATE 0 9.456e-17
C35 M1:GATE 0 4.931e-17
R36 M6:GATE M2:SRC 162.613 
R37 M2:SRC M7:SRC 74.6685 
CC29446 M2:SRC M12:GATE 5.75e-18
CC29464 M2:SRC M2:GATE 1.435e-17
CC29456 M2:SRC A2 6.848e-17
R38 M7:SRC M6:GATE 167.455 
CC29451 M7:SRC A2 1.185e-17
CC29439 M7:SRC M12:GATE 1.94e-17
R39 M6:GATE M9:GATE 139.125 
C40 M2:SRC 0 8.36e-18
C41 M7:SRC 0 7.94e-17
C42 M6:GATE 0 6.822e-17
C43 M9:GATE 0 3.413e-17
R44 A2 M12:GATE 152.373 
R45 M12:GATE M2:GATE 545.918 
R46 M2:GATE A2 118.665 
C47 M12:GATE 0 7.372e-17
C48 M2:GATE 0 5.748e-17
C49 A2 0 4.461e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
