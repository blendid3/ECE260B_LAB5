.SUBCKT MUX2D4 I0 I1 S Z
MMM20 M13:SRC M20:GATE M20:SRC vdd pch L=6e-08 W=4.15e-07  AD=4.8e-14  AS=5e-14  PD=7.98e-07  PS=6.7e-07  SA=6.62e-07  SB=2.26e-07  NRD=0.347  NRS=0.317  SCA=5.665  SCB=0.005  SCC=0.0001487 
MMM21 M20:SRC M21:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=6.4e-14  AS=5.2e-14  PD=8.5e-07  PS=7.2e-07  SA=4.25e-07  SB=3.74e-07  NRD=0.279  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 vdd M22:GATE M22:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.6e-14  PD=7.2e-07  PS=1.37e-06  SA=1.65e-07  SB=6.83e-07  NRD=2.099  NRS=0.433  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M9:SRC M10:GATE vss vss nch L=6e-08 W=3.9e-07  AD=4.4e-14  AS=3.9e-14  PD=7.14e-07  PS=5.9e-07  SA=4.25e-07  SB=3.25e-07  NRD=6.023  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.4e-14  PD=5.9e-07  PS=1.11e-06  SA=1.65e-07  SB=6.52e-07  NRD=4.183  NRS=0.575  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=5.4e-07  SB=1.16e-06  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vdd vdd pch L=6e-08 W=2.64e-07  AD=4.4e-14  AS=3.4e-14  PD=8.6e-07  PS=4.93e-07  SA=1.7e-07  SB=1.7e-06  NRD=0.737  NRS=0.658  SCA=15.255  SCB=0.017  SCC=0.002 
MMM2 M1:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=5.1e-14  PD=5.9e-07  PS=8.13e-07  SA=2.54e-07  SB=1.42e-06  NRD=4.183  NRS=5.397  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 M13:DRN M13:GATE M13:SRC vdd pch L=6e-08 W=3.43e-07  AD=5.6e-14  AS=4e-14  PD=1.01e-06  PS=6.62e-07  SA=3.38e-07  SB=1.65e-07  NRD=0.612  NRS=0.383  SCA=12.895  SCB=0.014  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=2.04e-07  AD=2.5e-14  AS=3.5e-14  PD=4.07e-07  PS=7.5e-07  SA=1.8e-07  SB=1.7e-06  NRD=0.797  NRS=0.972  SCA=18.109  SCB=0.02  SCC=0.002 
MMM14 M14:DRN M14:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=5.43e-07  SB=1.16e-06  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 vss M4:GATE M4:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=1.562e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 M14:DRN M15:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.8e-14  PD=7.2e-07  PS=9.87e-07  SA=2.58e-07  SB=1.42e-06  NRD=2.099  NRS=3.615  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 M5:DRN M5:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=1.299e-06  SB=4.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 vdd M16:GATE M16:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.562e-06  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 vss M6:GATE M6:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=1.056e-06  SB=6.6e-07  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 M17:DRN M17:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.3e-06  SB=4.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 M7:DRN M7:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=7.9e-07  SB=9.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 vdd M18:GATE M18:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=1.057e-06  SB=6.6e-07  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE M8:SRC vss nch L=6e-08 W=2.39e-07  AD=4.6e-14  AS=2.4e-14  PD=8.6e-07  PS=4.51e-07  SA=6.77e-07  SB=2e-07  NRD=1.436  NRS=0.768  SCA=5.844  SCB=0.005  SCC=9.292e-05 
MMM19 M19:DRN M19:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=7.92e-07  SB=9.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 M8:SRC M9:GATE M9:SRC vss nch L=6e-08 W=2.7e-07  AD=2.7e-14  AS=2.9e-14  PD=5.09e-07  PS=4.76e-07  SA=6.9e-07  SB=3.21e-07  NRD=6.681  NRS=0.46  SCA=6.917  SCB=0.007  SCC=0.000196 
R0 M16:SRC M17:DRN 0.001 
R1 M19:DRN M17:DRN 1301.35 
R2 M17:DRN Z 15.3562 
CC3990 M17:DRN M16:GATE 4.61e-17
CC3987 M17:DRN M17:GATE 4.509e-17
CC3972 M17:DRN N_12:1 1.102e-17
R3 M5:DRN Z 15.3454 
R4 M7:DRN Z 15.4574 
R5 Z M19:DRN 15.5392 
CC4009 Z M18:GATE 1.597e-17
CC4039 Z N_12:3 5.047e-17
CC4047 Z M7:GATE 1.161e-17
CC4002 Z M19:GATE 1.504e-17
CC3995 Z M4:GATE 7.64e-18
CC3992 Z M5:GATE 1.53e-17
CC3991 Z M16:GATE 6.35e-18
CC4052 Z M6:GATE 1.135e-17
CC3988 Z M17:GATE 2.094e-17
CC3982 Z N_12:2 4.91e-18
CC3977 Z N_12:1 4.667e-17
R6 M19:DRN M18:SRC 0.001 
CC4022 M19:DRN N_12:3 1.68e-18
CC4006 M19:DRN M18:GATE 4.6e-17
CC3998 M19:DRN M19:GATE 4.661e-17
CC3971 M19:DRN N_12:1 1.466e-17
R7 M6:SRC M7:DRN 0.001 
R8 M7:DRN M5:DRN 1337.66 
CC4032 M7:DRN N_12:3 1.678e-17
CC4044 M7:DRN M7:GATE 5.07e-18
CC4049 M7:DRN M6:GATE 6.77e-18
CC3975 M7:DRN N_12:1 8.83e-17
R9 M5:DRN M4:SRC 0.001 
CC4033 M5:DRN N_12:3 2.3e-18
CC3996 M5:DRN M4:GATE 8.48e-18
CC3993 M5:DRN M5:GATE 8.86e-18
CC3983 M5:DRN N_12:2 7.89e-17
CC3976 M5:DRN N_12:1 1.423e-17
C10 M17:DRN 0 1.361e-17
C11 Z 0 2.2992e-16
C12 M19:DRN 0 7.17e-18
C13 M7:DRN 0 5.21e-18
C14 M5:DRN 0 8.72e-18
R15 M3:SRC M13:GATE 379.453 
R16 M9:GATE M13:GATE 443.057 
R17 M13:GATE M12:DRN 379.817 
CC3880 M13:GATE M13:DRN 3.741e-17
CC3884 M13:GATE M8:DRN 3.29e-18
CC3890 M13:GATE M9:SRC 4.35e-18
CC3877 M13:GATE N_4:1 5.08e-18
CC4056 M13:GATE M8:SRC 1.146e-17
CC4013 M13:GATE M13:SRC 3.553e-17
CC4024 M13:GATE N_12:3 4.51e-18
CC3895 M13:GATE M20:GATE 4.95e-18
CC3904 M13:GATE M12:GATE 1.107e-17
CC3910 M13:GATE S 4.05e-18
CC3923 M13:GATE M8:GATE 3.11e-18
R18 M3:SRC M12:DRN 68.8761 
R19 M12:DRN M9:GATE 736.874 
CC3881 M12:DRN M13:DRN 1.204e-17
CC4026 M12:DRN N_12:3 2.916e-17
CC3878 M12:DRN N_4:1 4.051e-17
CC3906 M12:DRN M12:GATE 1.046e-17
CC3911 M12:DRN S 8.625e-17
R20 M9:GATE M3:SRC 736.159 
CC4029 M9:GATE N_12:3 2.107e-17
CC3888 M9:GATE M22:SRC 4.55e-18
CC3891 M9:GATE M9:SRC 3.015e-17
CC4058 M9:GATE M8:SRC 2.008e-17
CC3927 M9:GATE M8:GATE 2.13e-18
CC3882 M3:SRC M13:DRN 2.66e-18
CC3883 M3:SRC M8:DRN 1.725e-17
CC4061 M3:SRC M8:SRC 2.86e-18
CC4034 M3:SRC N_12:3 4.69e-18
CC3879 M3:SRC N_4:1 7.567e-17
CC4017 M3:SRC M13:SRC 5.06e-18
CC3899 M3:SRC M20:GATE 4.86e-18
CC3907 M3:SRC M12:GATE 2.1e-18
CC3919 M3:SRC M3:GATE 3.933e-17
CC3929 M3:SRC M8:GATE 7.45e-18
C21 M13:GATE 0 2.167e-17
C22 M12:DRN 0 1.019e-17
C23 M9:GATE 0 4.055e-17
C24 M3:SRC 0 1.008e-17
R25 N_4:1 M8:DRN 33.0596 
R26 M8:DRN M13:DRN 934.223 
CC3918 M8:DRN M3:GATE 1.376e-17
CC3928 M8:DRN M8:GATE 2.098e-17
CC4031 M8:DRN N_12:3 6.96e-18
R27 M13:DRN N_4:1 32.0922 
CC3905 M13:DRN M12:GATE 6.73e-18
CC3896 M13:DRN M20:GATE 1.7e-18
CC4025 M13:DRN N_12:3 5.37e-18
R28 M14:DRN N_4:1 30.1593 
R29 N_4:1 M1:DRN 31.4394 
CC3921 N_4:1 M3:GATE 2.37e-18
CC3915 N_4:1 S 8.14e-17
CC3908 N_4:1 M12:GATE 1.219e-17
CC3931 N_4:1 M8:GATE 3.29e-18
CC3954 N_4:1 I1:1 1.353e-17
CC3900 N_4:1 M20:GATE 3.83e-18
CC3959 N_4:1 M15:GATE 1.207e-17
CC3962 N_4:1 M14:GATE 5.3e-18
CC3967 N_4:1 I1 7.679e-17
CC3970 N_4:1 M2:GATE 5.6e-18
CC4018 N_4:1 M13:SRC 1.3e-18
CC4042 N_4:1 N_12:3 1.3059e-16
CC3952 M1:DRN I1:1 5.573e-17
CC3965 M1:DRN I1 1.641e-17
CC4038 M1:DRN N_12:3 1.426e-17
CC3947 M14:DRN I1:1 5.95e-18
CC3955 M14:DRN M15:GATE 2.865e-17
CC3960 M14:DRN M14:GATE 2.904e-17
CC3963 M14:DRN I1 2.91e-18
C30 M8:DRN 0 1.287e-17
C31 M13:DRN 0 9.63e-18
C32 N_4:1 0 1.0218e-16
C33 M14:DRN 0 5.95e-18
R34 M12:GATE S 110.333 
R35 S M3:GATE 94.962 
CC4040 S N_12:3 6.33e-18
CC3953 S I1:1 4.23e-18
CC3958 S M15:GATE 6.06e-18
CC3966 S I1 3.54e-18
R36 M12:GATE M3:GATE 270.952 
R37 M3:GATE M8:GATE 269.771 
CC3951 M3:GATE I1:1 6.93e-18
CC4035 M3:GATE N_12:3 6.93e-18
CC4059 M8:GATE M8:SRC 3.038e-17
CC3949 M8:GATE I1:1 7.97e-18
CC3969 M8:GATE M2:GATE 2.56e-18
CC4030 M8:GATE N_12:3 1.364e-17
R38 M12:GATE M20:GATE 416.052 
CC3957 M12:GATE M15:GATE 5.39e-18
CC3948 M12:GATE I1:1 5.95e-18
CC4015 M12:GATE M13:SRC 6.97e-18
CC3901 M12:GATE M22:SRC 5.22e-18
CC4012 M20:GATE M13:SRC 3.269e-17
CC4021 M20:GATE N_12:3 7.43e-18
CC3894 M20:GATE M20:SRC 3.869e-17
CC3893 M20:GATE M22:SRC 1.74e-18
C39 S 0 9.46e-18
C40 M3:GATE 0 3.045e-17
C41 M8:GATE 0 8.42e-17
C42 M12:GATE 0 1.0069e-16
C43 M20:GATE 0 5.851e-17
R44 M9:SRC M20:SRC 98.0627 
R45 M11:SRC M20:SRC 95.3922 
R46 M20:SRC M22:SRC 45.5755 
CC4020 M20:SRC N_12:3 3.968e-17
CC3939 M20:SRC M21:GATE 4.493e-17
CC3941 M20:SRC I0 8.995e-17
CC3933 M20:SRC I0:1 1.212e-17
R47 M9:SRC M22:SRC 94.1705 
R48 M22:SRC M11:SRC 91.606 
CC4053 M22:SRC M8:SRC 1.18e-18
CC4019 M22:SRC N_12:3 4.53e-18
CC3932 M22:SRC I0:1 2.41e-18
CC3944 M22:SRC M10:GATE 6.52e-18
CC3937 M22:SRC M22:GATE 6.199e-17
CC3938 M22:SRC M21:GATE 9.88e-18
CC3946 M22:SRC M11:GATE 7.26e-18
R49 M11:SRC M9:SRC 171.909 
CC4027 M11:SRC N_12:3 2.177e-17
CC3934 M11:SRC I0:1 2.795e-17
CC4028 M9:SRC N_12:3 1.06e-18
CC3945 M9:SRC M10:GATE 2.736e-17
CC3943 M9:SRC I0 1.35e-18
C50 M20:SRC 0 2.576e-17
C51 M22:SRC 0 1.1685e-16
C52 M11:SRC 0 6.236e-17
C53 M9:SRC 0 8.966e-17
R54 M22:GATE I0:1 111.3 
R55 M11:GATE I0:1 94.0755 
R56 I0 I0:1 38.5044 
R57 M10:GATE I0:1 203.073 
R58 I0:1 M21:GATE 240.255 
R59 I0 M21:GATE 436.522 
R60 M21:GATE M10:GATE 728.871 
R61 M10:GATE I0 368.964 
C62 I0:1 0 6.727e-17
C63 M21:GATE 0 6.591e-17
C64 M10:GATE 0 3.09e-17
C65 I0 0 3.169e-17
C66 M11:GATE 0 5.263e-17
C67 M22:GATE 0 5.864e-17
R68 M15:GATE I1:1 111.3 
R69 M2:GATE I1:1 94.0755 
R70 M14:GATE I1:1 270.681 
R71 M1:GATE I1:1 202.592 
R72 I1:1 I1 54.0381 
CC4043 I1:1 N_12:3 4.18e-18
CC3981 I1:1 N_12:1 6.28e-18
CC4048 I1:1 M7:GATE 6.19e-18
R73 M14:GATE I1 277.178 
R74 I1 M1:GATE 207.453 
CC4041 I1 N_12:3 4.026e-17
CC4003 I1 M19:GATE 2.06e-18
CC3979 I1 N_12:1 1.29e-18
R75 M1:GATE M14:GATE 1039.15 
CC4037 M1:GATE N_12:3 1.237e-17
CC4046 M1:GATE M7:GATE 4.02e-18
CC4000 M14:GATE M19:GATE 1.639e-17
CC4023 M14:GATE N_12:3 1.06e-18
CC3974 M14:GATE N_12:1 5.03e-18
CC4036 M2:GATE N_12:3 6.72e-18
C76 M15:GATE 0 5.258e-17
C77 I1:1 0 7.76e-18
C78 I1 0 1.88e-17
C79 M1:GATE 0 3.521e-17
C80 M14:GATE 0 4.146e-17
C81 M2:GATE 0 3.402e-17
R82 M8:SRC N_12:3 29.9999 
R83 M13:SRC N_12:3 30.8894 
R84 M7:GATE N_12:3 237.356 
R85 M19:GATE N_12:3 263.4 
R86 N_12:3 N_12:1 56.4615 
R87 M18:GATE N_12:1 84.8002 
R88 N_12:2 N_12:1 22.4472 
R89 M6:GATE N_12:1 98.0499 
R90 M7:GATE N_12:1 190.674 
R91 N_12:1 M19:GATE 211.593 
R92 M19:GATE M7:GATE 889.515 
R93 M5:GATE N_12:2 98.0499 
R94 M4:GATE N_12:2 144.585 
R95 M16:GATE N_12:2 158.261 
R96 N_12:2 M17:GATE 107.324 
R97 M16:GATE M4:GATE 638.114 
C98 M8:SRC 0 4.92e-18
C99 N_12:3 0 1.8186e-16
C100 N_12:1 0 1.769e-17
C101 M19:GATE 0 4.267e-17
C102 M7:GATE 0 2.923e-17
C103 M6:GATE 0 3.183e-17
C104 N_12:2 0 5.84e-18
C105 M17:GATE 0 3.757e-17
C106 M18:GATE 0 4.411e-17
C107 M13:SRC 0 1.22e-18
C108 M16:GATE 0 8.563e-17
C109 M4:GATE 0 5.925e-17
C110 M5:GATE 0 3.092e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
