.SUBCKT AN2D0 A1 A2 Z
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=1.95e-07  AD=3.9e-14  AS=1.6e-14  PD=7.9e-07  PS=3.55e-07  SA=2e-07  SB=7.6e-07  NRD=1.069  NRS=20.501  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM2 M1:SRC M2:GATE vss vss nch L=6e-08 W=1.98e-07  AD=1.6e-14  AS=2.9e-14  PD=3.55e-07  PS=4.95e-07  SA=4.2e-07  SB=5.4e-07  NRD=20.501  NRS=0.939  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM3 M3:DRN M3:GATE vss vss nch L=6e-08 W=2.02e-07  AD=3.5e-14  AS=2.9e-14  PD=7.5e-07  PS=4.95e-07  SA=7.8e-07  SB=1.8e-07  NRD=0.972  NRS=0.939  SCA=5.801  SCB=0.005  SCC=8.311e-05 
MMM4 vdd M4:GATE M4:SRC vdd pch L=6e-08 W=2.65e-07  AD=5.2e-14  AS=2.7e-14  PD=9.2e-07  PS=4.7e-07  SA=2e-07  SB=7.6e-07  NRD=0.84  NRS=0.438  SCA=6.553  SCB=0.007  SCC=0.00018 
MMM5 M4:SRC M5:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=2.7e-14  AS=3.2e-14  PD=4.7e-07  PS=5.1e-07  SA=4.7e-07  SB=4.9e-07  NRD=0.438  NRS=0.727  SCA=6.553  SCB=0.007  SCC=0.00018 
MMM6 M6:DRN M6:GATE vdd vdd pch L=6e-08 W=2.65e-07  AD=4.7e-14  AS=3.2e-14  PD=8.8e-07  PS=5.1e-07  SA=7.8e-07  SB=1.8e-07  NRD=0.771  NRS=0.727  SCA=6.553  SCB=0.007  SCC=0.00018 
R0 M3:DRN Z 30.4633 
R1 Z M6:DRN 30.488 
CC75162 Z M6:GATE 1.867e-17
CC75163 Z M4:SRC 8.71e-17
CC75164 Z M3:GATE 3.9e-18
CC75165 Z M1:DRN 1.22e-18
CC75166 M6:DRN M6:GATE 2.735e-17
CC75167 M6:DRN M4:SRC 1.61e-18
CC75169 M3:DRN M3:GATE 2.219e-17
CC75170 M3:DRN M4:SRC 8.17e-18
C2 Z 0 1.0527e-16
C3 M6:DRN 0 2.377e-17
C4 M3:DRN 0 2.09e-17
R5 M4:GATE M1:GATE 682.92 
R6 M1:GATE A1 155.757 
CC75158 M1:GATE M4:SRC 6.93e-18
CC75160 M1:GATE M2:GATE 4.82e-18
CC75161 M1:GATE M1:DRN 2.136e-17
R7 A1 M4:GATE 137.944 
CC75155 A1 M4:SRC 2.09e-18
CC75156 A1 M1:DRN 9.32e-18
CC75157 A1 A2 7.16e-17
CC75154 A1 M5:GATE 1.05e-18
CC75153 A1 M6:GATE 3.766e-17
CC75152 M4:GATE A2 6.52e-18
CC75150 M4:GATE M4:SRC 3.655e-17
CC75149 M4:GATE M5:GATE 8.62e-18
C8 M1:GATE 0 3.344e-17
C9 A1 0 4.701e-17
C10 M4:GATE 0 4.828e-17
R11 A2 M5:GATE 145.288 
R12 M5:GATE M2:GATE 666.771 
CC75140 M5:GATE M4:SRC 4.229e-17
CC75139 M5:GATE M6:GATE 7.48e-18
R13 M2:GATE A2 144.907 
CC75146 M2:GATE M4:SRC 1.649e-17
CC75145 M2:GATE M3:GATE 1.07e-18
CC75144 A2 M1:DRN 8.299e-17
CC75143 A2 M3:GATE 3.51e-18
CC75142 A2 M4:SRC 4.94e-18
CC75141 A2 M6:GATE 5.29e-18
C14 M5:GATE 0 3.642e-17
C15 M2:GATE 0 3.936e-17
C16 A2 0 1.893e-17
R17 M1:DRN M3:GATE 380.97 
R18 M4:SRC M3:GATE 374.987 
R19 M3:GATE M6:GATE 484.762 
R20 M1:DRN M6:GATE 337.401 
R21 M6:GATE M4:SRC 332.105 
R22 M4:SRC M1:DRN 75.7303 
C23 M3:GATE 0 7.567e-17
C24 M6:GATE 0 3.922e-17
C25 M4:SRC 0 5.101e-17
C26 M1:DRN 0 1.2674e-16
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
