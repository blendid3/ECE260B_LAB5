.SUBCKT BUFFD2 I Z
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.2e-14  AS=4.9e-14  PD=1.1e-06  PS=6.4e-07  SA=1.6e-07  SB=7.45e-07  NRD=0.567  NRS=0.654  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=6.8e-14  AS=3.9e-14  PD=1.13e-06  PS=5.9e-07  SA=7.3e-07  SB=1.75e-07  NRD=0.496  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=4.9e-14  AS=3.9e-14  PD=6.4e-07  PS=5.9e-07  SA=4.7e-07  SB=4.35e-07  NRD=0.654  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=8.3e-14  AS=6.5e-14  PD=1.36e-06  PS=7.7e-07  SA=1.6e-07  SB=7.45e-07  NRD=0.532  NRS=0.66  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vdd M5:GATE M5:SRC vdd pch L=6e-08 W=5.2e-07  AD=9.1e-14  AS=5.2e-14  PD=1.39e-06  PS=7.2e-07  SA=7.3e-07  SB=1.75e-07  NRD=0.446  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.5e-14  PD=7.2e-07  PS=7.7e-07  SA=4.7e-07  SB=4.35e-07  NRD=2.057  NRS=0.66  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M6:DRN Z 15.4602 
R1 Z M3:SRC 15.3048 
CC77792 Z M3:GATE 2.42e-18
CC77790 Z M1:DRN 1.748e-17
CC77771 Z N_8:1 2.696e-17
CC77774 Z M6:GATE 5.39e-18
CC77778 Z M5:GATE 7.45e-18
CC77782 Z M4:DRN 6.173e-17
CC77784 Z M2:GATE 3.92e-18
R2 M3:SRC M2:SRC 0.001 
CC77794 M3:SRC M3:GATE 8.11e-18
CC77788 M3:SRC M1:DRN 5.98e-18
CC77769 M3:SRC N_8:1 9.289e-17
CC77785 M3:SRC M2:GATE 8.55e-18
R3 M6:DRN M5:SRC 0.001 
CC77786 M6:DRN M1:DRN 1.82e-18
CC77768 M6:DRN N_8:1 1.66e-17
CC77775 M6:DRN M6:GATE 4.575e-17
CC77777 M6:DRN M5:GATE 4.576e-17
C4 Z 0 1.4811e-16
C5 M3:SRC 0 1.516e-17
C6 M6:DRN 0 7.94e-18
R7 M4:GATE M1:GATE 505.187 
R8 M1:GATE I 117.422 
CC77770 M1:GATE N_8:1 1.573e-17
CC77781 M1:GATE M4:DRN 2.71e-18
R9 I M4:GATE 143.544 
CC77772 I N_8:1 8.742e-17
CC77776 I M6:GATE 1.87e-18
CC77783 I M4:DRN 7.47e-18
CC77791 I M1:DRN 3.755e-17
CC77773 M4:GATE M6:GATE 4.76e-18
CC77780 M4:GATE M4:DRN 2.803e-17
CC77787 M4:GATE M1:DRN 1.136e-17
C10 M1:GATE 0 5.117e-17
C11 I 0 2.599e-17
C12 M4:GATE 0 7.713e-17
R13 M1:DRN M4:DRN 92.9663 
R14 M4:DRN N_8:1 92.9849 
R15 M3:GATE N_8:1 94.0755 
R16 M6:GATE N_8:1 111.3 
R17 M1:DRN N_8:1 92.4832 
R18 M5:GATE N_8:1 164.389 
R19 N_8:1 M2:GATE 138.947 
R20 M2:GATE M5:GATE 635.948 
C21 M4:DRN 0 7.782e-17
C22 N_8:1 0 2.841e-17
C23 M2:GATE 0 7.47e-17
C24 M5:GATE 0 1.0754e-16
C25 M1:DRN 0 9.885e-17
C26 M6:GATE 0 6.168e-17
C27 M3:GATE 0 5.598e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
