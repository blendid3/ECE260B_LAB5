.SUBCKT AN2D4 A1 A2 Z
MMM10 vdd M10:GATE M10:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.85e-07  SB=1.515e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM11 vdd M11:GATE M9:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.25e-07  SB=1.775e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.4e-14  AS=3.4e-14  PD=1.11e-06  PS=5.65e-07  SA=1.65e-07  SB=2.035e-06  NRD=0.575  NRS=7.952  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M10:SRC M12:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.45e-07  SB=1.255e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM2 M2:DRN M2:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.4e-14  PD=5.9e-07  PS=5.65e-07  SA=6.6e-07  SB=1.54e-06  NRD=4.183  NRS=7.952  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=2.04e-06  SB=1.6e-07  NRD=0.427  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 M2:DRN M3:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.4e-14  PD=5.9e-07  PS=5.65e-07  SA=4e-07  SB=1.8e-06  NRD=4.183  NRS=7.952  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=6.6e-14  PD=7.2e-07  PS=7.75e-07  SA=1.78e-06  SB=4.2e-07  NRD=2.099  NRS=0.315  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M2:SRC M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.4e-14  AS=4.9e-14  PD=5.65e-07  PS=6.4e-07  SA=8.95e-07  SB=1.305e-06  NRD=7.952  NRS=0.654  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vdd M15:GATE M15:SRC vdd pch L=6e-08 W=5.24e-07  AD=6.6e-14  AS=5.2e-14  PD=7.75e-07  PS=7.2e-07  SA=1.465e-06  SB=7.35e-07  NRD=0.315  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=2.04e-06  SB=1.6e-07  NRD=0.462  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.205e-06  SB=9.95e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=5e-14  PD=5.9e-07  PS=6.45e-07  SA=1.78e-06  SB=4.2e-07  NRD=4.183  NRS=0.654  SCA=11.955  SCB=0.013  SCC=0.001 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=5e-14  AS=3.9e-14  PD=6.45e-07  PS=5.9e-07  SA=1.465e-06  SB=7.35e-07  NRD=0.654  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=4.9e-14  PD=5.9e-07  PS=6.4e-07  SA=1.205e-06  SB=9.95e-07  NRD=4.183  NRS=0.654  SCA=11.955  SCB=0.013  SCC=0.001 
MMM9 vdd M9:GATE M9:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.6e-14  AS=5.2e-14  PD=1.37e-06  PS=7.2e-07  SA=1.65e-07  SB=2.035e-06  NRD=0.534  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 Z M5:SRC 30.2953 
R1 M5:SRC M6:DRN 0.001 
CC75719 M5:SRC N_11:2 5.634e-17
CC75712 M5:SRC N_11:1 1.315e-17
R2 Z M7:SRC 30.4161 
R3 M7:SRC M8:DRN 0.001 
CC75718 M7:SRC N_11:2 8.88e-18
CC75711 M7:SRC N_11:1 6.317e-17
R4 M13:SRC Z 30.4441 
R5 Z M15:SRC 30.5854 
CC75726 Z M16:GATE 2.14e-18
CC75744 Z M5:GATE 2.68e-18
CC75720 Z N_11:2 3.94e-18
CC75743 Z M6:GATE 8.31e-18
CC75715 Z N_11:1 1.1528e-16
CC75750 Z M2:DRN 5.21e-18
CC75746 Z M8:GATE 2.24e-18
CC75737 Z M13:GATE 6.64e-18
CC75735 Z M14:GATE 1.178e-17
CC75742 Z M7:GATE 7.63e-18
CC75731 Z M15:GATE 1.606e-17
R6 M15:SRC M16:DRN 0.001 
CC75724 M15:SRC M16:GATE 2.809e-17
CC75707 M15:SRC N_11:1 1.227e-17
CC75728 M15:SRC M15:GATE 2.797e-17
R7 M13:SRC M14:DRN 0.001 
CC75708 M13:SRC N_11:1 1.04e-17
CC75736 M13:SRC M13:GATE 2.806e-17
CC75734 M13:SRC M14:GATE 2.742e-17
C8 M5:SRC 0 6.09e-18
C9 M7:SRC 0 4.98e-18
C10 Z 0 1.8728e-16
C11 M15:SRC 0 7.28e-18
C12 M13:SRC 0 4.8e-18
R13 M12:GATE M4:GATE 506.173 
R14 M4:GATE A2:1 124.386 
CC75713 M4:GATE N_11:1 2.441e-17
CC75722 M4:GATE M10:SRC 1.15e-18
CC75784 M4:GATE M2:GATE 4.4e-18
CC75757 M4:GATE A1:1 9.21e-18
R15 M9:GATE A2:1 147.814 
R16 M1:GATE A2:1 113.551 
R17 A2 A2:1 0.2053 
R18 A2:1 M12:GATE 150.983 
CC75717 A2:1 N_11:1 2.799e-17
CC75764 A2:1 A1:1 3.078e-17
CC75776 A2:1 M10:GATE 1.109e-17
CC75740 A2:1 M9:SRC 2.069e-17
CC75783 A2:1 A1 7.898e-17
CC75751 A2:1 M2:DRN 9.067e-17
CC75727 A2:1 M16:GATE 2.07e-18
CC75723 A2:1 M10:SRC 3.93e-18
CC75788 A2:1 M3:GATE 5e-18
CC75709 M12:GATE N_11:1 7.57e-18
CC75721 M12:GATE M10:SRC 2.809e-17
CC75753 M12:GATE A1:1 4.04e-18
CC75773 M12:GATE M10:GATE 3.69e-18
CC75725 M12:GATE M16:GATE 6.76e-18
R19 M1:GATE M9:GATE 501.568 
CC75790 M1:GATE M3:GATE 5.11e-18
CC75761 M1:GATE A1:1 5.12e-18
CC75710 M9:GATE N_11:1 2.84e-18
CC75756 M9:GATE A1:1 1.018e-17
CC75738 M9:GATE M9:SRC 2.823e-17
CC75768 M9:GATE M11:GATE 7.94e-18
CC75780 M9:GATE A1 1.35e-18
C20 M4:GATE 0 3.21e-17
C21 A2:1 0 1.6292e-16
C22 M12:GATE 0 9.359e-17
C23 A2 0 3.9e-19
C24 M1:GATE 0 4.763e-17
C25 M9:GATE 0 7.921e-17
R26 N_11:2 M5:GATE 138.947 
R27 M5:GATE M13:GATE 635.948 
R28 M13:GATE N_11:2 164.389 
R29 M14:GATE N_11:2 111.3 
R30 N_11:1 N_11:2 63.4048 
R31 M7:GATE N_11:2 277.281 
R32 M15:GATE N_11:2 328.052 
R33 N_11:2 M6:GATE 94.0755 
R34 N_11:1 M15:GATE 239.529 
R35 M15:GATE M7:GATE 1047.51 
R36 M7:GATE N_11:1 202.458 
R37 M16:GATE N_11:1 111.3 
R38 M8:GATE N_11:1 82.8124 
R39 M10:SRC N_11:1 97.6312 
R40 M9:SRC N_11:1 100.22 
R41 N_11:1 M2:DRN 96.323 
CC75775 N_11:1 M10:GATE 5.29e-18
CC75763 N_11:1 A1:1 2.12e-18
CC75789 N_11:1 M3:GATE 2.11e-18
CC75770 N_11:1 M11:GATE 4.99e-18
CC75787 N_11:1 M2:GATE 3.62e-18
R42 M10:SRC M2:DRN 139.672 
R43 M2:DRN M9:SRC 143.375 
CC75792 M2:DRN M3:GATE 9.96e-18
CC75785 M2:DRN M2:GATE 2.97e-17
CC75760 M2:DRN A1:1 2.868e-17
R44 M9:SRC M10:SRC 127.204 
CC75755 M9:SRC A1:1 3.77e-18
CC75767 M9:SRC M11:GATE 2.79e-17
CC75779 M9:SRC A1 2.94e-18
CC75754 M10:SRC A1:1 3.126e-17
CC75778 M10:SRC A1 4.571e-17
C45 M5:GATE 0 7.06e-17
C46 M13:GATE 0 1.0652e-16
C47 N_11:2 0 2.987e-17
C48 M6:GATE 0 4.736e-17
C49 M15:GATE 0 7.451e-17
C50 M7:GATE 0 4.713e-17
C51 N_11:1 0 7.045e-17
C52 M2:DRN 0 4.404e-17
C53 M9:SRC 0 1.0421e-16
C54 M10:SRC 0 6.797e-17
C55 M8:GATE 0 2.063e-17
C56 M16:GATE 0 7.33e-17
C57 M14:GATE 0 7.32e-17
R58 M2:GATE M10:GATE 750.333 
R59 M10:GATE A1:1 155.07 
R60 M3:GATE A1:1 84.8002 
R61 M2:GATE A1:1 127.704 
R62 A1 A1:1 22 
R63 A1:1 M11:GATE 112.625 
C64 M10:GATE 0 6.113e-17
C65 A1:1 0 4.446e-17
C66 M11:GATE 0 6.859e-17
C67 A1 0 9.16e-18
C68 M2:GATE 0 2.984e-17
C69 M3:GATE 0 2.457e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
