.SUBCKT AN2D8 A1 A2 Z
MMM20 M18:SRC M20:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.44e-06  SB=2.16e-06  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 vdd M21:GATE M21:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=3.44e-06  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=3.18e-06  SB=4.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 vdd M23:GATE M23:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=2.94e-06  SB=6.6e-07  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 M24:DRN M24:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=2.68e-06  SB=9.2e-07  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM25 vdd M25:GATE M25:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=2.44e-06  SB=1.16e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM26 M26:DRN M26:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=2.18e-06  SB=1.42e-06  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM27 vdd M27:GATE M27:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=1.94e-06  SB=1.66e-06  NRD=6.61  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM28 M28:DRN M28:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=1.68e-06  SB=1.92e-06  NRD=2.057  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=2.68e-06  SB=9.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=2.44e-06  SB=1.16e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.6e-14  AS=2.9e-14  PD=1.12e-06  PS=5.4e-07  SA=1.7e-07  SB=3.43e-06  NRD=0.583  NRS=11.783  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=2.18e-06  SB=1.42e-06  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.97e-07  AD=5.3e-14  AS=2.9e-14  PD=6.6e-07  PS=5.4e-07  SA=7.1e-07  SB=2.89e-06  NRD=0.655  NRS=11.783  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vss M13:GATE M13:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=1.94e-06  SB=1.66e-06  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 vss M3:GATE M1:SRC vss nch L=6e-08 W=3.97e-07  AD=5.3e-14  AS=2.9e-14  PD=6.6e-07  PS=5.4e-07  SA=3.8e-07  SB=3.22e-06  NRD=0.655  NRS=11.783  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=4.5e-14  PD=5.9e-07  PS=6.2e-07  SA=1.68e-06  SB=1.92e-06  NRD=4.141  NRS=0.657  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 M4:DRN M4:GATE M4:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=2.9e-14  PD=5.9e-07  PS=5.4e-07  SA=1.18e-06  SB=2.42e-06  NRD=4.183  NRS=11.783  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vdd M15:GATE M15:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.6e-07  SB=3.44e-06  NRD=0.532  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 M4:DRN M5:GATE M2:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=2.9e-14  PD=5.9e-07  PS=5.4e-07  SA=9.2e-07  SB=2.68e-06  NRD=4.183  NRS=11.783  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 vdd M16:GATE M16:SRC vdd pch L=6e-08 W=5.24e-07  AD=4.7e-14  AS=5.2e-14  PD=7e-07  PS=7.2e-07  SA=6.6e-07  SB=2.94e-06  NRD=6.61  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M4:SRC M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=2.9e-14  AS=4.5e-14  PD=5.4e-07  PS=6.2e-07  SA=1.39e-06  SB=2.21e-06  NRD=11.783  NRS=0.657  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 M15:SRC M17:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=4.7e-14  PD=7.2e-07  PS=7e-07  SA=4.2e-07  SB=3.18e-06  NRD=2.099  NRS=6.61  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=3.44e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 vdd M18:GATE M18:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.18e-06  SB=2.42e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=3.18e-06  SB=4.2e-07  NRD=4.141  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vdd M19:GATE M16:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.2e-07  SB=2.68e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=2.94e-06  SB=6.6e-07  NRD=7.648  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
R0 M18:GATE M4:GATE 672.483 
R1 A1 M4:GATE 590.369 
R2 M4:GATE A1:1 185.518 
CC76365 M4:GATE M6:GATE 6.02e-18
CC76355 M4:GATE A2 1.762e-17
CC76375 M4:GATE N_21:3 5.88e-18
CC76420 M4:GATE M4:DRN 1.72e-18
R3 M5:GATE A1:1 98.0499 
R4 M18:GATE A1:1 203.068 
R5 A1 A1:1 33.9104 
R6 A1:1 M19:GATE 107.324 
CC76366 A1:1 M6:GATE 1.519e-17
CC76363 A1:1 M2:GATE 6.54e-18
CC76358 A1:1 A2 1.033e-17
CC76382 A1:1 N_21:3 6.9e-18
CC76349 A1:1 M16:GATE 4.64e-18
CC76340 A1:1 A2:1 2.51e-18
CC76425 A1:1 M4:DRN 5.495e-17
CC76368 M19:GATE N_21:3 4.41e-18
CC76345 M19:GATE M16:GATE 7.39e-18
CC76336 M19:GATE A2:1 1.33e-18
CC76394 M19:GATE M16:SRC 2.778e-17
R7 A1 M1:GATE 117.167 
R8 M1:GATE M15:GATE 502.788 
CC76359 M1:GATE M3:GATE 5.2e-18
CC76356 M1:GATE A2 4.69e-18
CC76378 M1:GATE N_21:3 6.08e-18
CC76338 M1:GATE A2:1 1.178e-17
CC76428 M1:GATE M1:DRN 6.13e-18
R9 M15:GATE A1 143.316 
CC76372 M15:GATE N_21:3 3.83e-18
CC76342 M15:GATE M17:GATE 7.48e-18
CC76337 M15:GATE A2:1 1.73e-18
CC76410 M15:GATE M15:SRC 2.811e-17
CC76426 M15:GATE M1:DRN 3.7e-18
R10 A1 M18:GATE 646.212 
CC76360 A1 M3:GATE 1.169e-17
CC76357 A1 A2 1.0795e-16
CC76380 A1 N_21:3 1.3255e-16
CC76348 A1 M16:GATE 5.98e-18
CC76343 A1 M17:GATE 7.76e-18
CC76339 A1 A2:1 1.069e-17
CC76423 A1 M4:DRN 7.24e-18
CC76399 A1 M16:SRC 7.38e-18
CC76429 A1 M1:DRN 2.902e-17
CC76413 A1 M15:SRC 7.62e-18
CC76369 M18:GATE N_21:3 7.21e-18
CC76353 M18:GATE A2 1.53e-18
CC76351 M18:GATE M20:GATE 7.52e-18
CC76389 M18:GATE M18:SRC 2.848e-17
CC76361 M5:GATE M2:GATE 1.701e-17
CC76374 M5:GATE N_21:3 1.03e-18
CC76419 M5:GATE M4:DRN 1.64e-18
C11 M4:GATE 0 2.472e-17
C12 A1:1 0 1.368e-17
C13 M19:GATE 0 8.543e-17
C14 M1:GATE 0 2.31e-17
C15 M15:GATE 0 7.293e-17
C16 A1 0 5.141e-17
C17 M18:GATE 0 7.717e-17
C18 M5:GATE 0 4.012e-17
R19 M20:GATE M6:GATE 519.657 
R20 M6:GATE A2 130.177 
CC76416 M6:GATE M14:GATE 7.71e-18
CC76373 M6:GATE N_21:3 8.96e-18
CC76390 M6:GATE M18:SRC 1.86e-18
R21 A2:1 A2 22.1342 
R22 A2 M20:GATE 144.352 
CC76405 A2 M28:GATE 1.74e-18
CC76422 A2 M4:DRN 6.21e-18
CC76412 A2 M15:SRC 1.15e-18
CC76391 A2 M18:SRC 4.6e-18
CC76379 A2 N_21:3 1.8393e-16
CC76367 M20:GATE N_21:3 1.368e-17
CC76383 M20:GATE N_21:4 6.67e-18
CC76387 M20:GATE M18:SRC 2.839e-17
CC76402 M20:GATE M28:GATE 1.541e-17
R23 M3:GATE A2:1 82.718 
CC76376 M3:GATE N_21:3 3.35e-18
R24 M17:GATE A2:1 111.3 
R25 M16:GATE A2:1 159.896 
R26 A2:1 M2:GATE 135.15 
CC76414 A2:1 M15:SRC 1.56e-18
CC76400 A2:1 M16:SRC 3.02e-18
CC76381 A2:1 N_21:3 4.5e-18
R27 M2:GATE M16:GATE 675.753 
CC76377 M2:GATE N_21:3 2.73e-18
CC76409 M16:GATE M15:SRC 1.04e-18
CC76371 M16:GATE N_21:3 1.43e-17
CC76397 M16:GATE M16:SRC 2.801e-17
CC76408 M17:GATE M15:SRC 2.79e-17
CC76370 M17:GATE N_21:3 6.99e-18
C28 M6:GATE 0 1.987e-17
C29 A2 0 4.055e-17
C30 M20:GATE 0 5.858e-17
C31 M3:GATE 0 2.637e-17
C32 A2:1 0 6.021e-17
C33 M2:GATE 0 3.889e-17
C34 M16:GATE 0 3.798e-17
C35 M17:GATE 0 3.674e-17
R36 M10:GATE N_21:1 98.0499 
R37 M24:GATE N_21:1 107.324 
R38 N_21:4 N_21:1 22.4472 
R39 M9:GATE N_21:1 250.804 
R40 M23:GATE N_21:1 274.53 
R41 N_21:1 N_21:2 57.4181 
CC76450 N_21:1 Z:1 8.21e-18
CC76487 N_21:1 M10:DRN 6.018e-17
R42 M22:GATE N_21:2 107.324 
R43 M8:GATE N_21:2 98.0499 
R44 M21:GATE N_21:2 158.261 
R45 M7:GATE N_21:2 144.585 
R46 M9:GATE N_21:2 231.512 
R47 N_21:2 M23:GATE 253.411 
CC76451 N_21:2 Z:1 4.5e-18
CC76488 N_21:2 M10:DRN 1.714e-17
CC76493 N_21:2 M8:DRN 7.556e-17
R48 M23:GATE M9:GATE 1106.92 
CC76459 M23:GATE Z:2 1.628e-17
CC76436 M23:GATE Z:1 5.89e-18
CC76475 M23:GATE M24:DRN 4.516e-17
CC76484 M9:GATE M10:DRN 1.266e-17
CC76443 M9:GATE Z:1 1.437e-17
R49 M14:GATE M28:GATE 893.526 
R50 N_21:3 M28:GATE 236.295 
R51 M28:GATE N_21:6 236.586 
CC76500 M28:GATE M28:DRN 4.61e-17
CC76454 M28:GATE Z:2 5.95e-18
CC76431 M28:GATE Z:1 2.32e-18
R52 M14:GATE N_21:6 213.354 
R53 M13:GATE N_21:6 87.8111 
R54 M27:GATE N_21:6 97.086 
R55 N_21:3 N_21:6 16.4019 
R56 N_21:6 N_21:5 21.5426 
CC76453 N_21:6 Z:1 5.2e-18
CC76523 N_21:6 M14:DRN 6.37e-17
R57 M26:GATE N_21:5 98.315 
R58 N_21:3 N_21:5 23.4332 
R59 M12:GATE N_21:5 89.0402 
R60 N_21:5 N_21:4 22.4472 
CC76452 N_21:5 Z:1 7.14e-18
CC76514 N_21:5 M12:DRN 4.256e-17
R61 M11:GATE N_21:4 98.0499 
R62 N_21:4 M25:GATE 84.8002 
CC76449 N_21:4 Z:1 4.911e-17
CC76467 N_21:4 Z:2 7.61e-18
CC76499 N_21:4 M26:DRN 1.272e-17
CC76481 N_21:4 M22:DRN 1.148e-17
CC76486 N_21:4 M10:DRN 1.529e-17
CC76492 N_21:4 M8:DRN 1.451e-17
CC76472 N_21:4 Z 1.062e-17
CC76477 N_21:4 M24:DRN 1.128e-17
CC76505 N_21:4 M28:DRN 1.267e-17
CC76512 N_21:4 M12:DRN 5.318e-17
CC76521 N_21:4 M14:DRN 1.423e-17
CC76457 M25:GATE Z:2 1.566e-17
CC76496 M25:GATE M26:DRN 4.518e-17
CC76434 M25:GATE Z:1 2.69e-18
CC76440 M12:GATE Z:1 1.1e-17
CC76508 M12:GATE M12:DRN 5.07e-18
R63 M14:GATE N_21:3 213.092 
R64 M4:DRN N_21:3 32.5225 
R65 M1:DRN N_21:3 33.9888 
R66 M15:SRC N_21:3 35.4057 
R67 M16:SRC N_21:3 34.6183 
R68 N_21:3 M18:SRC 33.0709 
CC76448 N_21:3 Z:1 9.768e-17
CC76471 N_21:3 Z 4.662e-17
CC76504 N_21:3 M28:DRN 2.15e-18
CC76520 N_21:3 M14:DRN 1.973e-17
R69 M15:SRC M18:SRC 999.39 
R70 M18:SRC M16:SRC 977.165 
CC76462 M18:SRC Z:2 7.9e-18
R71 M16:SRC M15:SRC 590.847 
CC76463 M16:SRC Z:2 6.32e-18
CC76464 M15:SRC Z:2 8.42e-18
CC76501 M27:GATE M28:DRN 4.497e-17
CC76455 M27:GATE Z:2 1.72e-17
R72 M1:DRN M4:DRN 791.054 
CC76447 M1:DRN Z:1 1.06e-18
CC76446 M4:DRN Z:1 7.65e-18
CC76456 M26:GATE Z:2 1.671e-17
CC76495 M26:GATE M26:DRN 4.53e-17
R73 M7:GATE M21:GATE 638.114 
CC76445 M7:GATE Z:1 5.51e-18
CC76491 M7:GATE M8:DRN 1.17e-17
CC76461 M21:GATE Z:2 5.96e-18
CC76480 M21:GATE M22:DRN 4.62e-17
CC76444 M8:GATE Z:1 1.575e-17
CC76490 M8:GATE M8:DRN 7.89e-18
CC76460 M22:GATE Z:2 1.894e-17
CC76479 M22:GATE M22:DRN 4.481e-17
CC76437 M22:GATE Z:1 1.76e-18
CC76441 M11:GATE Z:1 9.31e-18
CC76509 M11:GATE M12:DRN 9.19e-18
CC76458 M24:GATE Z:2 1.67e-17
CC76435 M24:GATE Z:1 3.96e-18
CC76474 M24:GATE M24:DRN 4.508e-17
CC76483 M10:GATE M10:DRN 5.01e-18
CC76442 M10:GATE Z:1 1.157e-17
CC76439 M13:GATE Z:1 1.098e-17
CC76518 M13:GATE M14:DRN 5.07e-18
CC76438 M14:GATE Z:1 2.12e-18
CC76517 M14:GATE M14:DRN 1.053e-17
C74 N_21:1 0 1.23e-18
C75 N_21:2 0 1.086e-17
C76 M23:GATE 0 2.893e-17
C77 M9:GATE 0 2.372e-17
C78 M28:GATE 0 3.52e-17
C79 N_21:6 0 1.88e-18
C80 N_21:5 0 1.74e-18
C81 N_21:4 0 5.463e-17
C82 M25:GATE 0 3.949e-17
C83 M12:GATE 0 3.147e-17
C84 N_21:3 0 2.4869e-16
C85 M18:SRC 0 7.54e-18
C86 M16:SRC 0 1.034e-17
C87 M15:SRC 0 1.722e-17
C88 M27:GATE 0 3.866e-17
C89 M1:DRN 0 1.456e-17
C90 M4:DRN 0 4.35e-18
C91 M26:GATE 0 4.039e-17
C92 M7:GATE 0 5.912e-17
C93 M21:GATE 0 7.788e-17
C94 M8:GATE 0 3.221e-17
C95 M22:GATE 0 2.387e-17
C96 M11:GATE 0 3.121e-17
C97 M24:GATE 0 5.184e-17
C98 M10:GATE 0 4.086e-17
C99 M13:GATE 0 3.084e-17
C100 M14:GATE 0 2.303e-17
R101 Z:1 Z 0.17333 
R102 Z:2 Z 0.25252 
R103 M26:DRN Z 53.5031 
R104 Z M28:DRN 52.2808 
R105 Z:2 M28:DRN 21.669 
R106 M28:DRN M27:SRC 0.001 
R107 Z:2 M26:DRN 21.4251 
R108 M26:DRN M25:SRC 0.001 
R109 Z:1 M14:DRN 15.2186 
R110 M14:DRN M13:SRC 0.001 
R111 M22:DRN Z:2 15.1709 
R112 Z:2 M24:DRN 14.9999 
R113 M24:DRN M23:SRC 0.001 
R114 M22:DRN M21:SRC 0.001 
R115 M10:DRN Z:1 15.0408 
R116 M8:DRN Z:1 15.1914 
R117 Z:1 M12:DRN 15.095 
R118 M12:DRN M11:SRC 0.001 
R119 M8:DRN M7:SRC 0.001 
R120 M10:DRN M9:SRC 0.001 
C121 Z 0 5.971e-17
C122 M28:DRN 0 4.84e-18
C123 M26:DRN 0 4.81e-18
C124 M14:DRN 0 1.96e-18
C125 Z:2 0 1.5393e-16
C126 M24:DRN 0 8.5e-18
C127 M22:DRN 0 1.026e-17
C128 Z:1 0 2.1108e-16
C129 M12:DRN 0 1.96e-18
C130 M8:DRN 0 2.91e-18
C131 M10:DRN 0 2.4e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
