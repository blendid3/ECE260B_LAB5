.SUBCKT AN2XD1 A1 A2 Z
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=7.8e-14  AS=3.1e-14  PD=1.18e-06  PS=5.5e-07  SA=2e-07  SB=7.6e-07  NRD=0.638  NRS=10.251  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M1:SRC M2:GATE vss vss nch L=6e-08 W=3.93e-07  AD=3.1e-14  AS=5.8e-14  PD=5.5e-07  PS=6.9e-07  SA=4.2e-07  SB=5.4e-07  NRD=10.251  NRS=0.662  SCA=11.955  SCB=0.013  SCC=0.001 
MMM3 M3:DRN M3:GATE vss vss nch L=6e-08 W=3.97e-07  AD=7e-14  AS=5.8e-14  PD=1.14e-06  PS=6.9e-07  SA=7.8e-07  SB=1.8e-07  NRD=0.6  NRS=0.662  SCA=11.955  SCB=0.013  SCC=0.001 
MMM4 vdd M4:GATE M4:SRC vdd pch L=6e-08 W=5.24e-07  AD=1.04e-13  AS=5.5e-14  PD=1.44e-06  PS=7.3e-07  SA=2e-07  SB=7.6e-07  NRD=0.564  NRS=0.287  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 M4:SRC M5:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.5e-14  AS=6.5e-14  PD=7.3e-07  PS=7.7e-07  SA=4.7e-07  SB=4.9e-07  NRD=0.287  NRS=0.66  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=9.4e-14  AS=6.5e-14  PD=1.4e-06  PS=7.7e-07  SA=7.8e-07  SB=1.8e-07  NRD=0.453  NRS=0.66  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 M6:DRN Z 15.4371 
CC9230 M6:DRN M6:GATE 4.578e-17
CC9222 M6:DRN M4:SRC 2.63e-18
R1 Z M3:DRN 30.4633 
CC9233 Z M6:GATE 1.252e-17
CC9240 Z M1:DRN 8.77e-17
CC9238 Z M3:GATE 5.75e-18
CC9225 M3:DRN M4:SRC 2.202e-17
CC9236 M3:DRN M3:GATE 6.68e-18
C2 M6:DRN 0 3.232e-17
C3 Z 0 1.0389e-16
C4 M3:DRN 0 2.608e-17
R5 A1 M4:GATE 142.288 
R6 M4:GATE M1:GATE 538.172 
CC9215 M4:GATE M5:GATE 6.49e-18
CC9224 M4:GATE M4:SRC 2.944e-17
CC9216 M4:GATE A2 1.41e-18
R7 M1:GATE A1 124.451 
CC9227 M1:GATE M4:SRC 9.69e-18
CC9220 M1:GATE M2:GATE 5.03e-18
CC9221 M1:GATE A2 1.544e-17
CC9242 A1 M1:DRN 3.263e-17
CC9229 A1 M4:SRC 2.08e-18
CC9235 A1 M6:GATE 3.227e-17
CC9217 A1 M5:GATE 5.64e-18
CC9218 A1 M2:GATE 1.004e-17
CC9219 A1 A2 4.423e-17
C8 M4:GATE 0 9.089e-17
C9 M1:GATE 0 2.901e-17
C10 A1 0 3.718e-17
R11 M1:DRN M6:GATE 352.267 
R12 M3:GATE M6:GATE 389.273 
R13 M6:GATE M4:SRC 350.034 
CC9231 M6:GATE M5:GATE 5.21e-18
R14 M1:DRN M4:SRC 76.653 
R15 M4:SRC M3:GATE 306.158 
CC9228 M4:SRC A2 1.766e-17
CC9223 M4:SRC M5:GATE 4.639e-17
CC9226 M4:SRC M2:GATE 1.95e-17
R16 M3:GATE M1:DRN 308.111 
CC9239 M3:GATE A2 1.441e-17
CC9241 M1:DRN A2 5.853e-17
C17 M6:GATE 0 6.673e-17
C18 M4:SRC 0 8.854e-17
C19 M3:GATE 0 8.091e-17
C20 M1:DRN 0 5.362e-17
R21 M5:GATE M2:GATE 516.931 
R22 M2:GATE A2 113.833 
R23 A2 M5:GATE 151.109 
C24 M2:GATE 0 2.833e-17
C25 A2 0 4.6e-17
C26 M5:GATE 0 6.618e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
