.SUBCKT ND2D1 A1 A2 ZN
MMM1 M1:DRN M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.6e-14  AS=3.9e-14  PD=1.12e-06  PS=5.9e-07  SA=4.3e-07  SB=1.7e-07  NRD=0.583  NRS=4.12  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM2 vss M2:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.6e-14  AS=3.9e-14  PD=1.12e-06  PS=5.9e-07  SA=1.7e-07  SB=4.3e-07  NRD=0.583  NRS=4.12  SCA=10.357  SCB=0.011  SCC=0.0008048 
MMM3 vdd M3:GATE M3:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.8e-14  AS=5.2e-14  PD=1.38e-06  PS=7.2e-07  SA=4.3e-07  SB=1.7e-07  NRD=0.538  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 vdd M4:GATE M4:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.8e-14  AS=5.2e-14  PD=1.38e-06  PS=7.2e-07  SA=1.7e-07  SB=4.3e-07  NRD=0.538  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
R0 A1 M1:GATE 118.894 
R1 M1:GATE M3:GATE 552.68 
CC44940 M1:GATE M1:DRN 8.81e-18
CC44947 M1:GATE A2 1.026e-17
CC44953 M1:GATE M2:GATE 3.47e-18
CC44939 M1:GATE ZN 1.567e-17
R2 M3:GATE A1 152.48 
CC44942 M3:GATE M4:GATE 2.16e-18
CC44946 M3:GATE A2 1.206e-17
CC44934 M3:GATE M4:SRC 5.12e-17
CC44935 M3:GATE ZN 7.68e-18
CC44950 A1 A2 1.459e-17
CC44951 A1 M2:GATE 6.97e-18
CC44937 A1 M1:DRN 2.355e-17
CC44938 A1 ZN 7.724e-17
CC44936 A1 M4:SRC 1.102e-17
C3 M1:GATE 0 2.136e-17
C4 M3:GATE 0 8.296e-17
C5 A1 0 4.016e-17
R6 M4:GATE M2:GATE 531.535 
R7 M2:GATE A2 120.181 
CC44952 M2:GATE ZN 1.86e-18
R8 A2 M4:GATE 146.033 
CC44945 A2 M4:SRC 5.97e-18
CC44949 A2 ZN 1.707e-17
CC44941 M4:GATE M4:SRC 5.139e-17
CC44943 M4:GATE ZN 4.49e-18
C9 M2:GATE 0 4.969e-17
C10 A2 0 1.0116e-16
C11 M4:GATE 0 9.416e-17
R12 ZN M4:SRC 15.923 
R13 M4:SRC M3:SRC 0.001 
R14 ZN M1:DRN 30.5301 
C15 M4:SRC 0 1.979e-17
C16 ZN 0 1.6553e-16
C17 M1:DRN 0 2.644e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
