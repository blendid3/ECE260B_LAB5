.SUBCKT INVD12 I ZN
MMM20 M20:DRN M20:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.225e-06  SB=1.96e-06  NRD=2.099  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 vdd M21:GATE M21:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.6e-07  SB=2.24e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=7e-07  SB=2.5e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 vdd M23:GATE M23:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.4e-07  SB=2.76e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 M24:DRN M24:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=9.4e-14  PD=7.2e-07  PS=1.4e-06  SA=1.8e-07  SB=3.02e-06  NRD=2.057  NRS=0.545  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M10:DRN M10:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=7e-07  SB=2.5e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 vss M11:GATE M11:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.4e-07  SB=2.76e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=3.9e-07  AD=6.2e-14  AS=3.9e-14  PD=1.1e-06  PS=5.9e-07  SA=3.04e-06  SB=1.6e-07  NRD=0.462  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M12:DRN M12:GATE vss vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=7e-14  PD=5.9e-07  PS=1.14e-06  SA=1.8e-07  SB=3.02e-06  NRD=4.141  NRS=0.6  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 M2:DRN M2:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.78e-06  SB=4.2e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=3.04e-06  SB=1.6e-07  NRD=0.427  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 vss M3:GATE M3:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.52e-06  SB=6.8e-07  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.78e-06  SB=4.2e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2.26e-06  SB=9.4e-07  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vdd M15:GATE M15:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.52e-06  SB=6.8e-07  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 vss M5:GATE M5:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=2e-06  SB=1.2e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2.26e-06  SB=9.4e-07  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M6:DRN M6:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.74e-06  SB=1.46e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 vdd M17:GATE M17:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=2e-06  SB=1.2e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 vss M7:GATE M7:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.48e-06  SB=1.72e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M18:DRN M18:GATE vdd vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.74e-06  SB=1.46e-06  NRD=2.057  NRS=2.534  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M8:DRN M8:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.22e-06  SB=1.98e-06  NRD=4.141  NRS=4.537  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vdd M19:GATE M19:SRC vdd pch L=6e-08 W=5.24e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.48e-06  SB=1.72e-06  NRD=2.534  NRS=2.057  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 vss M9:GATE M9:SRC vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.6e-07  SB=2.24e-06  NRD=4.537  NRS=4.141  SCA=11.955  SCB=0.013  SCC=0.001 
R0 M23:GATE I:11 101.061 
CC9317 M23:GATE M24:DRN 4.519e-17
CC9245 M23:GATE ZN:1 1.586e-17
R1 I I:11 70.5223 
R2 I:10 I:11 21.5119 
R3 M11:GATE I:11 83.8364 
R4 I:6 I:11 32.4825 
R5 I:11 I:2 22.3616 
CC9357 I:11 M12:DRN 4.082e-17
R6 I I:2 35.0797 
R7 M12:GATE I:2 80.5597 
R8 M24:GATE I:2 97.7846 
R9 I:2 I:6 60.8432 
CC9355 I:2 M12:DRN 2.54e-17
R10 I I:6 0.73013 
R11 I:5 I:6 40.1243 
R12 I:10 I:6 22 
R13 I:6 I:7 18.1946 
CC9368 I:6 M10:DRN 1.35e-18
CC9292 I:6 ZN:2 9.581e-17
CC9321 I:6 M24:DRN 1.57e-18
CC9329 I:6 M22:DRN 1.55e-18
CC9264 I:6 ZN:1 8.271e-17
CC9359 I:6 M12:DRN 1.16e-18
R14 M9:GATE I:7 82.8124 
R15 I:5 I:7 33.618 
R16 I:10 I:7 21.9794 
R17 I:7 M21:GATE 100.037 
CC9369 I:7 M10:DRN 4.067e-17
CC9326 M21:GATE M22:DRN 4.495e-17
CC9247 M21:GATE ZN:1 1.7e-17
R18 M1:GATE I:3 94.0755 
CC9286 M1:GATE ZN:2 2.06e-18
CC9307 M1:GATE M2:DRN 4.8e-18
R19 M13:GATE I:3 111.3 
R20 I:8 I:3 213.181 
R21 I:9 I:3 167.713 
R22 I:3 I:1 27.1529 
CC9310 I:3 M2:DRN 4.114e-17
CC9298 I:3 ZN:2 2.85e-18
R23 I:8 I:1 85.1358 
R24 M2:GATE I:1 94.0755 
R25 I:9 I:1 23.0504 
R26 I:1 M14:GATE 111.3 
CC9337 I:1 M20:DRN 4.99e-18
CC9309 I:1 M2:DRN 3.777e-17
CC9322 I:1 M24:DRN 2.63e-18
CC9297 I:1 ZN:2 1.78e-18
CC9330 I:1 M22:DRN 4.88e-18
CC9269 I:1 ZN:1 2.758e-17
CC9301 M14:GATE M14:DRN 4.479e-17
CC9254 M14:GATE ZN:1 1.755e-17
CC9316 M24:GATE M24:DRN 4.606e-17
CC9244 M24:GATE ZN:1 4.15e-18
CC9276 M11:GATE ZN:2 1.376e-17
CC9352 M11:GATE M12:DRN 4.59e-18
R27 M15:GATE I:9 88.7752 
R28 I:8 I:9 16.5354 
R29 I:9 M3:GATE 81.9458 
CC9365 I:9 M10:DRN 1.643e-17
CC9289 I:9 ZN:2 1.0526e-16
CC9335 I:9 M20:DRN 1.112e-17
CC9347 I:9 M4:DRN 5.855e-17
CC9342 I:9 M18:DRN 1.111e-17
CC9320 I:9 M24:DRN 1.105e-17
CC9308 I:9 M2:DRN 1.761e-17
CC9303 I:9 M14:DRN 1.247e-17
CC9315 I:9 M16:DRN 1.266e-17
CC9328 I:9 M22:DRN 1.114e-17
CC9261 I:9 ZN:1 6.715e-17
CC9356 I:9 M12:DRN 1.614e-17
CC9386 I:9 M6:DRN 1.631e-17
CC9376 I:9 M8:DRN 1.64e-17
CC9345 M3:GATE M4:DRN 4.57e-18
CC9284 M3:GATE ZN:2 6.35e-18
R30 M22:GATE I:10 103.792 
R31 I:10 M10:GATE 86.5669 
CC9367 I:10 M10:DRN 4.077e-17
CC9291 I:10 ZN:2 1.26e-18
CC9277 M10:GATE ZN:2 1.563e-17
CC9361 M10:GATE M10:DRN 4.57e-18
CC9275 M12:GATE ZN:2 3.76e-18
CC9351 M12:GATE M12:DRN 2.095e-17
CC9285 M2:GATE ZN:2 1.273e-17
CC9306 M2:GATE M2:DRN 7.33e-18
R32 M6:GATE I:4 94.0755 
CC9281 M6:GATE ZN:2 1.191e-17
CC9383 M6:GATE M6:DRN 4.57e-18
R33 M18:GATE I:4 111.3 
R34 M17:GATE I:4 282.501 
R35 M19:GATE I:4 275.689 
R36 I:8 I:4 58.1624 
R37 M5:GATE I:4 238.78 
R38 I:5 I:4 60.2341 
R39 I:4 M7:GATE 233.022 
CC9295 I:4 ZN:2 2.78e-18
CC9267 I:4 ZN:1 4.47e-18
CC9387 I:4 M6:DRN 5.943e-17
CC9381 I:4 M8:DRN 1.987e-17
R40 M19:GATE M7:GATE 1066.52 
R41 M7:GATE I:5 233.022 
CC9373 M7:GATE M8:DRN 4.57e-18
CC9280 M7:GATE ZN:2 1.303e-17
CC9256 M7:GATE ZN:1 1.28e-18
R42 M20:GATE I:5 111.3 
R43 M19:GATE I:5 275.689 
R44 I:5 M8:GATE 94.0755 
CC9266 I:5 ZN:1 2.06e-18
CC9380 I:5 M8:DRN 6.255e-17
CC9372 M8:GATE M8:DRN 4.57e-18
CC9279 M8:GATE ZN:2 1.566e-17
R45 M17:GATE M5:GATE 1092.88 
R46 M5:GATE I:8 225.005 
CC9282 M5:GATE ZN:2 1.16e-17
CC9258 M5:GATE ZN:1 1.65e-18
CC9384 M5:GATE M6:DRN 5.38e-18
R47 M16:GATE I:8 103.792 
R48 M17:GATE I:8 266.204 
R49 I:8 M4:GATE 86.5669 
CC9348 I:8 M4:DRN 4.06e-17
CC9296 I:8 ZN:2 3.071e-17
CC9268 I:8 ZN:1 3.725e-17
CC9388 I:8 M6:DRN 2.186e-17
CC9344 M4:GATE M4:DRN 4.49e-18
CC9283 M4:GATE ZN:2 8.55e-18
CC9362 M9:GATE M10:DRN 4.57e-18
CC9278 M9:GATE ZN:2 1.406e-17
CC9287 I ZN:2 2.33e-18
CC9259 I ZN:1 4.98e-18
CC9333 M19:GATE M20:DRN 4.485e-17
CC9249 M19:GATE ZN:1 2.451e-17
CC9340 M17:GATE M18:DRN 4.507e-17
CC9274 M17:GATE ZN:2 2.63e-18
CC9251 M17:GATE ZN:1 1.752e-17
CC9312 M16:GATE M16:DRN 4.476e-17
CC9252 M16:GATE ZN:1 1.776e-17
CC9313 M15:GATE M16:DRN 4.499e-17
CC9253 M15:GATE ZN:1 1.797e-17
CC9325 M22:GATE M22:DRN 4.557e-17
CC9246 M22:GATE ZN:1 1.859e-17
CC9302 M13:GATE M14:DRN 4.597e-17
CC9255 M13:GATE ZN:1 5.15e-18
CC9339 M18:GATE M18:DRN 4.478e-17
CC9250 M18:GATE ZN:1 2.235e-17
CC9332 M20:GATE M20:DRN 4.538e-17
CC9248 M20:GATE ZN:1 1.835e-17
C50 M23:GATE 0 4.001e-17
C51 I:11 0 4.14e-18
C52 I:2 0 3.519e-17
C53 I:6 0 1.449e-17
C54 I:7 0 1.237e-17
C55 M21:GATE 0 4.6e-17
C56 M1:GATE 0 5.853e-17
C57 I:3 0 2.736e-17
C58 I:1 0 1.85e-17
C59 M14:GATE 0 1.581e-17
C60 M24:GATE 0 6.508e-17
C61 M11:GATE 0 3.155e-17
C62 I:9 0 1.1644e-16
C63 M3:GATE 0 3.828e-17
C64 I:10 0 9.52e-18
C65 M10:GATE 0 3.211e-17
C66 M12:GATE 0 2.588e-17
C67 M2:GATE 0 3.271e-17
C68 M6:GATE 0 3.233e-17
C69 I:4 0 2.73e-18
C70 M7:GATE 0 3.968e-17
C71 I:5 0 5.23e-18
C72 M8:GATE 0 2.899e-17
C73 M5:GATE 0 3.093e-17
C74 I:8 0 2.93e-18
C75 M4:GATE 0 3.317e-17
C76 M9:GATE 0 2.557e-17
C77 I 0 7.034e-17
C78 M19:GATE 0 5.121e-17
C79 M17:GATE 0 4.376e-17
C80 M16:GATE 0 4.571e-17
C81 M15:GATE 0 4.667e-17
C82 M22:GATE 0 5.113e-17
C83 M13:GATE 0 5.747e-17
C84 M18:GATE 0 4.529e-17
C85 M20:GATE 0 4.489e-17
R86 ZN:2 M8:DRN 15.3688 
R87 M8:DRN M7:SRC 0.001 
R88 ZN:1 M18:DRN 14.9999 
R89 M18:DRN M17:SRC 0.001 
R90 M12:DRN M10:DRN 763.182 
R91 ZN:2 M10:DRN 15.6177 
R92 M10:DRN M9:SRC 0.001 
R93 ZN:1 M20:DRN 15.3575 
R94 M20:DRN M19:SRC 0.001 
R95 M23:SRC M24:DRN 0.001 
R96 ZN:1 M24:DRN 15.7864 
R97 M24:DRN M22:DRN 786.479 
R98 ZN:1 M22:DRN 15.5985 
R99 M22:DRN M21:SRC 0.001 
R100 M16:DRN ZN:1 15.4762 
R101 M14:DRN ZN:1 15.6625 
R102 ZN:1 ZN 0.104 
R103 ZN ZN:2 0.03813 
R104 M12:DRN ZN:2 15.8118 
R105 M6:DRN ZN:2 14.9999 
R106 M4:DRN ZN:2 15.4916 
R107 ZN:2 M2:DRN 15.6841 
R108 M4:DRN M2:DRN 951.315 
R109 M2:DRN M1:SRC 0.001 
R110 M4:DRN M3:SRC 0.001 
R111 M13:SRC M14:DRN 0.001 
R112 M14:DRN M16:DRN 980.689 
R113 M16:DRN M15:SRC 0.001 
R114 M5:SRC M6:DRN 0.001 
R115 M11:SRC M12:DRN 0.001 
C116 M8:DRN 0 1.95e-18
C117 M18:DRN 0 4.32e-18
C118 M10:DRN 0 2e-18
C119 M20:DRN 0 4.32e-18
C120 M24:DRN 0 2.78e-17
C121 M22:DRN 0 1.189e-17
C122 ZN:1 0 3.0079e-16
C123 ZN 0 2.3e-19
C124 ZN:2 0 2.8944e-16
C125 M2:DRN 0 3.76e-18
C126 M4:DRN 0 2.17e-18
C127 M14:DRN 0 1.096e-17
C128 M16:DRN 0 4e-18
C129 M6:DRN 0 1.9e-18
C130 M12:DRN 0 4.93e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
