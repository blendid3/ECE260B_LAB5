.SUBCKT OAI21D4 A1 A2 B ZN
MMM20 M19:SRC M20:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=7.4e-14  PD=7.2e-07  PS=1.39e-06  SA=1.39e-07  SB=1.98e-06  NRD=2.099  NRS=0.525  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM21 M21:DRN M21:GATE M21:SRC vdd pch L=6e-08 W=5.2e-07  AD=7.7e-14  AS=5.2e-14  PD=1.37e-06  PS=7.2e-07  SA=9.4e-07  SB=1.47e-07  NRD=0.527  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM22 M22:DRN M22:GATE M22:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.8e-07  SB=4.08e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM23 M22:SRC M23:GATE M23:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.2e-07  SB=6.68e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM24 M24:DRN M24:GATE M24:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=8.3e-14  PD=7.2e-07  PS=1.36e-06  SA=1.6e-07  SB=9.28e-07  NRD=2.099  NRS=0.427  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM10 M9:SRC M10:GATE M10:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=6.8e-07  SB=1.465e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM11 M11:DRN M11:GATE M11:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=4.2e-07  SB=1.725e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM1 M1:DRN M1:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.2e-14  AS=3.5e-14  PD=1.1e-06  PS=5.7e-07  SA=9.05e-07  SB=1.6e-07  NRD=0.567  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM12 M11:SRC M12:GATE M12:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=6.2e-14  PD=5.9e-07  PS=1.1e-06  SA=1.6e-07  SB=1.985e-06  NRD=4.183  NRS=0.567  SCA=11.955  SCB=0.013  SCC=0.001 
MMM2 vss M2:GATE M2:SRC vss nch L=6e-08 W=3.97e-07  AD=3.5e-14  AS=3.9e-14  PD=5.7e-07  PS=5.9e-07  SA=6.65e-07  SB=4e-07  NRD=7.648  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM13 vdd M13:GATE M13:SRC vdd pch L=6e-08 W=5.2e-07  AD=8.3e-14  AS=5.2e-14  PD=1.36e-06  PS=7.2e-07  SA=1.962e-06  SB=1.6e-07  NRD=0.532  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM3 M2:SRC M3:GATE vss vss nch L=6e-08 W=3.97e-07  AD=3.9e-14  AS=3.5e-14  PD=5.9e-07  PS=5.7e-07  SA=4.05e-07  SB=6.6e-07  NRD=4.183  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM14 M14:DRN M14:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.702e-06  SB=4.2e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM4 M4:DRN M4:GATE vss vss nch L=6e-08 W=3.97e-07  AD=6.4e-14  AS=3.5e-14  PD=1.11e-06  PS=5.7e-07  SA=1.65e-07  SB=9e-07  NRD=0.575  NRS=7.648  SCA=11.955  SCB=0.013  SCC=0.001 
MMM15 vdd M15:GATE M15:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.442e-06  SB=6.8e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM5 M5:DRN M5:GATE M5:SRC vss nch L=6e-08 W=3.9e-07  AD=6.4e-14  AS=3.9e-14  PD=1.11e-06  PS=5.9e-07  SA=1.98e-06  SB=1.65e-07  NRD=0.575  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM16 M16:DRN M16:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=1.182e-06  SB=9.4e-07  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM6 M5:SRC M6:GATE M6:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.72e-06  SB=4.25e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM17 vdd M17:GATE M17:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=9.22e-07  SB=1.2e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM7 M7:DRN M7:GATE M7:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.46e-06  SB=6.85e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM18 M17:SRC M18:GATE vdd vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=6.62e-07  SB=1.46e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM8 M7:SRC M8:GATE M8:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=1.2e-06  SB=9.45e-07  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
MMM19 vdd M19:GATE M19:SRC vdd pch L=6e-08 W=5.2e-07  AD=5.2e-14  AS=5.2e-14  PD=7.2e-07  PS=7.2e-07  SA=4.01e-07  SB=1.72e-06  NRD=2.099  NRS=2.099  SCA=9.643  SCB=0.01  SCC=0.000823 
MMM9 M9:DRN M9:GATE M9:SRC vss nch L=6e-08 W=3.9e-07  AD=3.9e-14  AS=3.9e-14  PD=5.9e-07  PS=5.9e-07  SA=9.4e-07  SB=1.205e-06  NRD=4.183  NRS=4.183  SCA=11.955  SCB=0.013  SCC=0.001 
R0 M14:GATE B:2 111.3 
CC92927 M14:GATE ZN:2 7.13e-18
CC92934 M14:GATE M13:SRC 2.17e-18
R1 M2:GATE B:2 86.5669 
R2 B B:2 22 
R3 B:1 B:2 21.4183 
R4 M1:GATE B:2 135.84 
R5 B:2 M13:GATE 160.712 
CC92998 B:2 M2:SRC 2.046e-17
CC92932 B:2 ZN:2 1.41e-18
CC92938 B:2 M13:SRC 2.594e-17
CC93029 B:2 M1:DRN 1.796e-17
R6 M13:GATE M1:GATE 667.973 
CC92928 M13:GATE ZN:2 5.23e-18
CC92935 M13:GATE M13:SRC 2.832e-17
CC93014 M1:GATE N_36:2 9.01e-18
CC93026 M1:GATE M1:DRN 1.152e-17
R7 M15:GATE B:1 111.3 
CC92926 M15:GATE ZN:2 4.41e-18
R8 M3:GATE B:1 81.5607 
R9 M4:GATE B:1 137.629 
R10 M16:GATE B:1 143.632 
R11 B:1 B 22.1714 
CC92943 B:1 M5:DRN 2.67e-18
CC92997 B:1 M2:SRC 2.832e-17
CC92937 B:1 M13:SRC 5.42e-18
CC92941 B:1 M15:SRC 4.422e-17
CC93064 B:1 M4:DRN 2.292e-17
CC93022 B:1 N_36:2 9.72e-18
CC92995 B M2:SRC 1.73e-18
CC92930 B ZN:2 4.166e-17
CC93016 B N_36:2 2.104e-17
R12 M16:GATE M4:GATE 455.169 
CC92925 M16:GATE ZN:2 1.223e-17
CC92933 M16:GATE M13:SRC 4.19e-18
CC92939 M16:GATE M15:SRC 2.787e-17
CC92929 M4:GATE ZN:2 2.704e-17
CC93061 M4:GATE M4:DRN 9.18e-18
CC93011 M4:GATE N_36:2 1.33e-18
CC92993 M2:GATE M2:SRC 9.13e-18
CC93013 M2:GATE N_36:2 8.18e-18
CC92992 M3:GATE M2:SRC 9.13e-18
CC93012 M3:GATE N_36:2 8.3e-18
C13 M14:GATE 0 3.91e-17
C14 B:2 0 2.694e-17
C15 M13:GATE 0 5.742e-17
C16 M1:GATE 0 3.474e-17
C17 M15:GATE 0 5.597e-17
C18 B:1 0 5.138e-17
C19 B 0 2.223e-17
C20 M16:GATE 0 1.0539e-16
C21 M4:GATE 0 4.954e-17
C22 M2:GATE 0 2.016e-17
C23 M3:GATE 0 2.261e-17
R24 M11:DRN M10:SRC 0.001 
R25 M10:SRC ZN:1 29.9999 
CC93005 M10:SRC N_36:2 5.69e-18
CC92953 M10:SRC A1:2 2.935e-17
CC92947 M10:SRC A1:1 1.865e-17
CC92979 M10:SRC M11:GATE 2.413e-17
R26 M12:SRC ZN:1 30.325 
R27 M6:SRC ZN:1 102.355 
R28 ZN ZN:1 0.11281 
R29 M8:SRC ZN:1 49.7221 
R30 ZN:1 ZN:2 2.62089 
CC93037 ZN:1 M11:SRC 1.53e-18
CC92956 ZN:1 A1:2 1.76e-18
CC92964 ZN:1 M23:GATE 1.512e-17
CC92960 ZN:1 M24:GATE 3.57e-18
CC92950 ZN:1 A1:1 2.878e-17
CC93152 ZN:1 M22:SRC 2.83e-18
CC92980 ZN:1 M11:GATE 4.17e-18
CC92985 ZN:1 M9:GATE 1.14e-18
CC93138 ZN:1 N_11:1 1.592e-17
CC92968 ZN:1 M22:GATE 1.65e-18
CC92977 ZN:1 A1 1.82e-17
R31 M13:SRC ZN:2 33.4092 
R32 M15:SRC ZN:2 32.5906 
R33 M6:SRC ZN:2 44.1278 
R34 M5:DRN ZN:2 29.9999 
R35 ZN:2 M8:SRC 79.5565 
CC93039 ZN:2 M11:SRC 6.44e-18
CC93021 ZN:2 N_36:2 2.6192e-16
CC93092 ZN:2 A2:3 4.13e-18
CC93081 ZN:2 M17:GATE 1.426e-17
CC93116 ZN:2 M7:GATE 2.31e-18
CC93117 ZN:2 M8:GATE 3.11e-18
CC93102 ZN:2 M6:GATE 2.31e-18
CC93101 ZN:2 A2 9.285e-17
CC93058 ZN:2 M5:SRC 5.95e-18
CC93055 ZN:2 M7:SRC 5.97e-18
CC93050 ZN:2 M9:SRC 5.97e-18
CC93063 ZN:2 M4:DRN 7.8e-18
CC93161 ZN:2 M24:SRC 9.55e-18
CC93188 ZN:2 M17:SRC 1.31e-17
CC93183 ZN:2 M19:SRC 4.89e-18
CC92951 ZN:2 A1:1 1.141e-17
CC92982 ZN:2 M10:GATE 2.31e-18
CC92972 ZN:2 M21:GATE 2.69e-18
CC92978 ZN:2 A1 4.265e-17
R36 M8:SRC M9:DRN 0.001 
CC93008 M8:SRC N_36:2 5.69e-18
CC93071 M8:SRC A2:2 3.026e-17
CC92983 M8:SRC M9:GATE 2.525e-17
CC92975 M8:SRC A1 6.18e-18
CC93010 M5:DRN N_36:2 5.84e-18
CC93087 M5:DRN A2:3 1.37e-17
CC93080 M5:DRN M17:GATE 4.53e-18
CC93107 M5:DRN M5:GATE 2.484e-17
CC93097 M5:DRN A2 2.86e-18
CC93060 M5:DRN M4:DRN 7.69e-18
R37 M24:DRN M23:SRC 0.001 
R38 M23:SRC ZN 30.3575 
CC92958 M23:SRC M24:GATE 2.791e-17
CC92961 M23:SRC M23:GATE 2.75e-17
CC93122 M23:SRC N_11:1 5.65e-18
CC93154 M23:SRC M24:SRC 1e-18
CC92944 M23:SRC A1:1 8.56e-18
R39 ZN M21:SRC 30.7688 
CC92959 ZN M24:GATE 1.71e-18
CC92967 ZN M22:GATE 3.87e-18
CC92963 ZN M23:GATE 3.47e-18
CC92949 ZN A1:1 6.42e-18
CC93149 ZN M22:SRC 6.14e-18
CC93134 ZN N_11:1 1.0864e-16
CC92970 ZN M21:GATE 1.82e-18
CC92976 ZN A1 9.85e-18
R40 M21:SRC M22:DRN 0.001 
CC92966 M21:SRC M22:GATE 2.823e-17
CC92945 M21:SRC A1:1 8.87e-18
CC92969 M21:SRC M21:GATE 2.821e-17
CC93125 M21:SRC N_11:1 5.9e-18
R41 M7:DRN M6:SRC 0.001 
CC93009 M6:SRC N_36:2 5.69e-18
CC93085 M6:SRC A2:3 1.121e-17
CC93078 M6:SRC M17:GATE 3.76e-18
CC93112 M6:SRC M7:GATE 4.66e-18
CC93095 M6:SRC A2 3.61e-18
CC93073 M6:SRC A2:2 2.519e-17
CC93066 M6:SRC A2:1 2.937e-17
CC93156 M12:SRC M24:SRC 1.51e-18
CC92946 M12:SRC A1:1 2.954e-17
CC93131 M12:SRC N_11:1 1.44e-18
R42 M13:SRC M15:SRC 764.335 
R43 M15:SRC M16:DRN 0.001 
R44 M13:SRC M14:DRN 0.001 
C45 M10:SRC 0 1.56e-18
C46 ZN:1 0 1.184e-17
C47 ZN:2 0 1.1343e-16
C48 M8:SRC 0 1.92e-18
C49 M5:DRN 0 4.54e-18
C50 M23:SRC 0 3.42e-18
C51 ZN 0 7.77e-18
C52 M21:SRC 0 1.069e-17
C53 M6:SRC 0 1.91e-18
C54 M12:SRC 0 7.7e-18
C55 M15:SRC 0 2.048e-17
C56 M13:SRC 0 2.295e-17
R57 M24:GATE A1:1 111.3 
CC93121 M24:GATE N_11:1 9.22e-18
CC93153 M24:GATE M24:SRC 4.378e-17
R58 M12:GATE A1:1 94.0755 
R59 A1:2 A1:1 60.2341 
R60 M11:GATE A1:1 233.022 
R61 A1:1 M23:GATE 275.689 
CC93137 A1:1 N_11:1 2.59e-18
CC93151 A1:1 M22:SRC 1.119e-17
CC93158 A1:1 M24:SRC 3.7e-18
CC93018 A1:1 N_36:2 2.21e-18
CC93036 A1:1 M11:SRC 9.63e-18
CC93047 A1:1 M9:SRC 7.18e-18
R62 A1:2 M23:GATE 275.689 
R63 M23:GATE M11:GATE 1066.52 
CC93144 M23:GATE M22:SRC 2.931e-17
CC93123 M23:GATE N_11:1 5.91e-18
R64 M11:GATE A1:2 233.022 
CC93033 M11:GATE M11:SRC 9.46e-18
CC93004 M11:GATE N_36:2 5.54e-18
R65 M10:GATE A1:2 94.0755 
R66 M22:GATE A1:2 111.3 
R67 A1 A1:2 37.0768 
R68 M9:GATE A1:2 199.267 
R69 A1:2 M21:GATE 235.753 
CC93172 A1:2 M21:DRN 4.41e-18
CC93038 A1:2 M11:SRC 1.764e-17
CC93049 A1:2 M9:SRC 1.891e-17
R70 A1 M21:GATE 462.113 
R71 M21:GATE M9:GATE 715.482 
CC93126 M21:GATE N_11:1 1.127e-17
CC93164 M21:GATE M21:DRN 2.479e-17
R72 M9:GATE A1 390.595 
CC93044 M9:GATE M9:SRC 9.46e-18
CC93007 M9:GATE N_36:2 5.54e-18
CC93136 A1 N_11:1 2.06e-17
CC93170 A1 M21:DRN 1.08e-18
CC93017 A1 N_36:2 2.83e-18
CC93046 A1 M9:SRC 2.25e-18
CC93145 M22:GATE M22:SRC 2.938e-17
CC93124 M22:GATE N_11:1 6.03e-18
CC93043 M10:GATE M9:SRC 2.962e-17
CC93006 M10:GATE N_36:2 6.18e-18
CC93032 M12:GATE M11:SRC 3.022e-17
CC93003 M12:GATE N_36:2 4.44e-18
C73 M24:GATE 0 2.903e-17
C74 A1:1 0 2.508e-17
C75 M23:GATE 0 2.585e-17
C76 M11:GATE 0 1.577e-17
C77 A1:2 0 8.22e-18
C78 M21:GATE 0 5.021e-17
C79 M9:GATE 0 2.849e-17
C80 A1 0 2.208e-17
C81 M22:GATE 0 3.424e-17
C82 M10:GATE 0 2.192e-17
C83 M12:GATE 0 2.304e-17
R84 N_36:1 M7:SRC 45.8448 
R85 M7:SRC N_36:2 92.724 
CC93084 M7:SRC A2:3 7.06e-18
CC93111 M7:SRC M7:GATE 9.46e-18
CC93120 M7:SRC M8:GATE 2.962e-17
CC93077 M7:SRC M17:GATE 1.77e-18
CC93072 M7:SRC A2:2 2.019e-17
R86 M11:SRC N_36:2 29.9999 
R87 N_36:1 N_36:2 2.09325 
R88 N_36:2 M9:SRC 45.3387 
CC93089 N_36:2 A2:3 5.03e-18
CC93103 N_36:2 M6:GATE 6.08e-18
CC93099 N_36:2 A2 5.44e-18
CC93109 N_36:2 M5:GATE 1.61e-18
CC93118 N_36:2 M8:GATE 6.32e-18
CC93114 N_36:2 M7:GATE 5.3e-18
R89 M9:SRC N_36:1 92.724 
R90 M5:SRC N_36:1 29.9999 
R91 M4:DRN N_36:1 31.9622 
R92 M2:SRC N_36:1 33.3351 
R93 N_36:1 M1:DRN 34.0586 
R94 M4:DRN M1:DRN 1508.68 
R95 M1:DRN M2:SRC 760.713 
R96 M2:SRC M4:DRN 1476.62 
CC93088 M4:DRN A2:3 1.21e-18
CC93108 M4:DRN M5:GATE 1.32e-18
CC93086 M5:SRC A2:3 2.507e-17
CC93105 M5:SRC M6:GATE 2.982e-17
CC93106 M5:SRC M5:GATE 9.54e-18
CC93079 M5:SRC M17:GATE 3.42e-18
C97 M7:SRC 0 5.4e-18
C98 N_36:2 0 2.7527e-16
C99 M9:SRC 0 1.2e-17
C100 N_36:1 0 1.175e-17
C101 M1:DRN 0 1.407e-17
C102 M2:SRC 0 4.1e-19
C103 M4:DRN 0 1.071e-17
C104 M5:SRC 0 5.4e-18
C105 M11:SRC 0 5.93e-18
R106 M5:GATE A2:3 85.7767 
R107 A2:1 A2:3 32.9458 
R108 M17:GATE A2:3 129.257 
R109 A2 A2:3 17.2395 
R110 A2:3 M18:GATE 111.3 
CC93187 A2:3 M17:SRC 6.639e-17
CC93141 A2:3 N_11:1 1.489e-17
CC93182 A2:3 M19:SRC 9.73e-18
CC93175 A2:3 M21:DRN 3e-18
CC93129 M18:GATE N_11:1 6.48e-18
R111 A2:1 A2 22.0421 
R112 A2 A2:2 17.4789 
CC93135 A2 N_11:1 5.588e-17
CC93185 A2 M17:SRC 1.26e-18
R113 M8:GATE A2:2 114.84 
R114 M20:GATE A2:2 111.3 
R115 A2:1 A2:2 32.7038 
R116 A2:2 M7:GATE 81.5607 
R117 M19:GATE A2:1 111.3 
R118 A2:1 M6:GATE 94.0755 
CC93140 A2:1 N_11:1 1.98e-18
CC93181 A2:1 M19:SRC 2.789e-17
CC93165 M20:GATE M21:DRN 3.1e-18
CC93177 M20:GATE M19:SRC 2.814e-17
CC93127 M20:GATE N_11:1 8.95e-18
CC93128 M19:GATE N_11:1 5.1e-18
C119 M5:GATE 0 1.809e-17
C120 A2:3 0 9.626e-17
C121 M18:GATE 0 5.241e-17
C122 A2 0 2.514e-17
C123 A2:2 0 1.388e-17
C124 M7:GATE 0 2.959e-17
C125 M17:GATE 0 5.487e-17
C126 A2:1 0 3.541e-17
C127 M6:GATE 0 2.372e-17
C128 M20:GATE 0 7.357e-17
C129 M19:GATE 0 5.874e-17
C130 M8:GATE 0 2.696e-17
R131 M22:SRC N_11:1 29.9999 
R132 M24:SRC N_11:1 15.8083 
R133 M19:SRC N_11:1 35.7175 
R134 M21:DRN N_11:1 33.5348 
R135 N_11:1 M17:SRC 36.6269 
R136 M19:SRC M17:SRC 484.52 
R137 M17:SRC M21:DRN 887.347 
R138 M21:DRN M19:SRC 865.317 
C139 N_11:1 0 2.2228e-16
C140 M17:SRC 0 4.6e-18
C141 M21:DRN 0 1.38e-17
C142 M19:SRC 0 1.387e-17
C143 M24:SRC 0 2.15e-17
C144 M22:SRC 0 8.27e-18
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
