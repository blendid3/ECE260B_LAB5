.SUBCKT NR2D0 A1 A2 ZN
MMM1 vss M1:GATE M1:SRC vss nch L=6e-08 W=1.95e-07  AD=3.6e-14  AS=2e-14  PD=7.6e-07  PS=3.95e-07  SA=4.45e-07  SB=1.85e-07  NRD=0.996  NRS=8.262  SCA=5.69  SCB=0.005  SCC=7.614e-05 
MMM2 vss M2:GATE M1:SRC vss nch L=6e-08 W=1.95e-07  AD=3.6e-14  AS=2e-14  PD=7.6e-07  PS=3.95e-07  SA=1.85e-07  SB=4.45e-07  NRD=0.996  NRS=8.262  SCA=5.69  SCB=0.005  SCC=7.614e-05 
MMM3 M3:DRN M3:GATE M3:SRC vdd pch L=6e-08 W=2.6e-07  AD=4.4e-14  AS=2.6e-14  PD=8.6e-07  PS=4.6e-07  SA=4.3e-07  SB=1.7e-07  NRD=0.737  NRS=4.018  SCA=4.967  SCB=0.004  SCC=5.833e-05 
MMM4 vdd M4:GATE M3:SRC vdd pch L=6e-08 W=2.6e-07  AD=4.4e-14  AS=2.6e-14  PD=8.6e-07  PS=4.6e-07  SA=1.7e-07  SB=4.3e-07  NRD=0.737  NRS=4.018  SCA=4.967  SCB=0.004  SCC=5.833e-05 
R0 M3:DRN ZN 30.5557 
R1 ZN M1:SRC 30.8956 
CC47584 ZN M1:GATE 2.06e-18
CC47582 ZN A1 8.97e-17
CC47592 ZN A2 1.84e-17
CC47579 ZN M3:GATE 9.48e-18
CC47590 M1:SRC A2 8.54e-18
CC47583 M1:SRC M1:GATE 2.3e-17
CC47581 M1:SRC A1 1.088e-17
CC47594 M1:SRC M2:GATE 2.307e-17
CC47577 M3:DRN M3:GATE 3.037e-17
C2 ZN 0 1.4636e-16
C3 M1:SRC 0 9.61e-18
C4 M3:DRN 0 2.386e-17
R5 M1:GATE A1 150.589 
R6 A1 M3:GATE 162.756 
CC47593 A1 A2 2.268e-17
CC47597 A1 M2:GATE 6.72e-18
CC47588 A1 M4:GATE 1.312e-17
R7 M3:GATE M1:GATE 800.708 
CC47589 M3:GATE A2 3.9e-18
CC47585 M3:GATE M4:GATE 1.134e-17
CC47591 M1:GATE A2 1.266e-17
CC47595 M1:GATE M2:GATE 2.01e-18
C8 A1 0 3.609e-17
C9 M3:GATE 0 4.36e-17
C10 M1:GATE 0 4.248e-17
R11 A2 M2:GATE 146.757 
R12 M2:GATE M4:GATE 755.135 
R13 M4:GATE A2 159.043 
C14 M2:GATE 0 4.859e-17
C15 M4:GATE 0 7.62e-17
C16 A2 0 9.638e-17
.ENDS
*.SCALE METER
.GLOBAL VSS VDD
